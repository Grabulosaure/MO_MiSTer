LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
PACKAGE rom_pack IS

  TYPE arr8  IS ARRAY(natural RANGE<>) OF unsigned(7 DOWNTO 0);

  CONSTANT ROM_BASIC6_0 : arr8 := (
    x"D5",x"D9",x"D6",x"08",x"D5",x"9E",x"CA",x"6A",x"D6",x"AB",x"D6",x"F1",x"D7",x"34",x"D7",x"AE",
    x"D7",x"B5",x"D8",x"0B",x"CC",x"D4",x"CC",x"11",x"CB",x"64",x"CB",x"9F",x"CC",x"0E",x"CC",x"5B",
    x"E3",x"BE",x"D6",x"27",x"21",x"E9",x"21",x"F9",x"D5",x"E0",x"22",x"3C",x"21",x"F9",x"E8",x"9F",
    x"E8",x"B1",x"CC",x"52",x"CC",x"25",x"CC",x"1E",x"CC",x"67",x"CC",x"E7",x"D0",x"D9",x"DB",x"B6",
    x"E4",x"6E",x"E3",x"DE",x"E4",x"69",x"E7",x"14",x"E7",x"1B",x"E4",x"36",x"E8",x"AD",x"22",x"DB",
    x"26",x"EB",x"28",x"23",x"2E",x"EB",x"C1",x"D4",x"C2",x"D0",x"C5",x"19",x"C7",x"E5",x"C8",x"00",
    x"FF",x"AE",x"04",x"00",x"00",x"03",x"02",x"79",x"D2",x"AC",x"79",x"D2",x"9F",x"7C",x"D2",x"EE",
    x"7C",x"D5",x"1C",x"7F",x"D6",x"B4",x"50",x"C8",x"86",x"46",x"C8",x"8C",x"3C",x"C8",x"92",x"32",
    x"C8",x"9D",x"28",x"C8",x"98",x"7A",x"D3",x"77",x"7B",x"D3",x"4A",x"64",x"C8",x"7F",x"64",x"C8",
    x"65",x"64",x"C8",x"6D",x"D3",x"D4",x"C8",x"79",x"D5",x"D4",x"C8",x"73",x"D5",x"D3",x"C8",x"7C",
    x"45",x"4E",x"C4",x"46",x"4F",x"D2",x"4E",x"45",x"58",x"D4",x"44",x"41",x"54",x"C1",x"44",x"49",
    x"CD",x"52",x"45",x"41",x"C4",x"FF",x"47",x"CF",x"52",x"55",x"CE",x"49",x"C6",x"52",x"45",x"53",
    x"54",x"4F",x"52",x"C5",x"52",x"45",x"54",x"55",x"52",x"CE",x"52",x"45",x"CD",x"A7",x"53",x"54",
    x"4F",x"D0",x"45",x"4C",x"53",x"C5",x"54",x"52",x"4F",x"CE",x"54",x"52",x"4F",x"46",x"C6",x"44",
    x"45",x"46",x"53",x"54",x"D2",x"44",x"45",x"46",x"49",x"4E",x"D4",x"44",x"45",x"46",x"53",x"4E",
    x"C7",x"FF",x"4F",x"CE",x"54",x"55",x"4E",x"C5",x"45",x"52",x"52",x"4F",x"D2",x"52",x"45",x"53",
    x"55",x"4D",x"C5",x"41",x"55",x"54",x"CF",x"44",x"45",x"4C",x"45",x"54",x"C5",x"4C",x"4F",x"43",
    x"41",x"54",x"C5",x"43",x"4C",x"D3",x"43",x"4F",x"4E",x"53",x"4F",x"4C",x"C5",x"50",x"53",x"45",
    x"D4",x"4D",x"4F",x"54",x"4F",x"D2",x"53",x"4B",x"49",x"50",x"C6",x"45",x"58",x"45",x"C3",x"42",
    x"45",x"45",x"D0",x"43",x"4F",x"4C",x"4F",x"D2",x"4C",x"49",x"4E",x"C5",x"42",x"4F",x"D8",x"FF",
    x"41",x"54",x"54",x"52",x"C2",x"44",x"45",x"C6",x"50",x"4F",x"4B",x"C5",x"50",x"52",x"49",x"4E",
    x"D4",x"43",x"4F",x"4E",x"D4",x"4C",x"49",x"53",x"D4",x"43",x"4C",x"45",x"41",x"D2",x"44",x"4F",
    x"D3",x"FF",x"4E",x"45",x"D7",x"53",x"41",x"56",x"C5",x"4C",x"4F",x"41",x"C4",x"4D",x"45",x"52",
    x"47",x"C5",x"4F",x"50",x"45",x"CE",x"43",x"4C",x"4F",x"53",x"C5",x"49",x"4E",x"50",x"45",x"CE",
    x"50",x"45",x"CE",x"50",x"4C",x"41",x"D9",x"54",x"41",x"42",x"A8",x"54",x"CF",x"53",x"55",x"C2",
    x"46",x"CE",x"53",x"50",x"43",x"A8",x"55",x"53",x"49",x"4E",x"C7",x"55",x"53",x"D2",x"45",x"52",
    x"CC",x"45",x"52",x"D2",x"4F",x"46",x"C6",x"54",x"48",x"45",x"CE",x"4E",x"4F",x"D4",x"53",x"54",
    x"45",x"D0",x"AB",x"AD",x"AA",x"AF",x"DE",x"41",x"4E",x"C4",x"4F",x"D2",x"58",x"4F",x"D2",x"45",
    x"51",x"D6",x"49",x"4D",x"D0",x"4D",x"4F",x"C4",x"C0",x"BE",x"BD",x"BC",x"53",x"47",x"CE",x"49",
    x"4E",x"D4",x"41",x"42",x"D3",x"46",x"52",x"C5",x"53",x"51",x"D2",x"4C",x"4F",x"C7",x"45",x"58",
    x"D0",x"43",x"4F",x"D3",x"53",x"49",x"CE",x"54",x"41",x"CE",x"50",x"45",x"45",x"CB",x"4C",x"45",
    x"CE",x"53",x"54",x"52",x"A4",x"56",x"41",x"CC",x"41",x"53",x"C3",x"43",x"48",x"52",x"A4",x"45",
    x"4F",x"C6",x"43",x"49",x"4E",x"D4",x"FF",x"FF",x"46",x"49",x"D8",x"48",x"45",x"58",x"A4",x"FF",
    x"53",x"54",x"49",x"43",x"CB",x"53",x"54",x"52",x"49",x"C7",x"47",x"52",x"A4",x"4C",x"45",x"46",
    x"54",x"A4",x"52",x"49",x"47",x"48",x"54",x"A4",x"4D",x"49",x"44",x"A4",x"49",x"4E",x"53",x"54",
    x"D2",x"56",x"41",x"52",x"50",x"54",x"D2",x"52",x"4E",x"C4",x"49",x"4E",x"4B",x"45",x"59",x"A4",
    x"49",x"4E",x"50",x"55",x"D4",x"43",x"53",x"52",x"4C",x"49",x"CE",x"50",x"4F",x"49",x"4E",x"D4",
    x"53",x"43",x"52",x"45",x"45",x"CE",x"50",x"4F",x"D3",x"50",x"54",x"52",x"49",x"C7",x"00",x"C4",
    x"9E",x"CF",x"97",x"D0",x"5C",x"C5",x"E2",x"CA",x"61",x"DD",x"3B",x"21",x"F9",x"C5",x"5F",x"C5",
    x"4B",x"C5",x"EA",x"C4",x"8A",x"C5",x"C1",x"C5",x"E5",x"C5",x"E5",x"C4",x"A7",x"C5",x"E5",x"CF",
    x"1F",x"CF",x"20",x"CE",x"EC",x"CE",x"EF",x"CE",x"E9",x"21",x"F9",x"C6",x"1F",x"F4",x"F3",x"CF",
    x"24",x"CF",x"2D",x"22",x"36",x"CE",x"C5",x"E5",x"FE",x"E8",x"FC",x"E6",x"40",x"E7",x"93",x"EC",
    x"6C",x"EB",x"CE",x"E8",x"E9",x"E8",x"FA",x"E6",x"B3",x"E8",x"1B",x"E8",x"2C",x"21",x"F9",x"E6",
    x"1C",x"E8",x"68",x"CC",x"DD",x"CD",x"7A",x"C4",x"CF",x"E0",x"6A",x"C4",x"DE",x"F1",x"94",x"21",
    x"F9",x"C4",x"22",x"E0",x"A3",x"E2",x"8C",x"E2",x"58",x"E1",x"E9",x"E1",x"B8",x"E8",x"C3",x"21",
    x"F9",x"EF",x"28",x"4F",x"4B",x"0D",x"0A",x"00",x"0D",x"0A",x"42",x"72",x"65",x"61",x"6B",x"00",
    x"45",x"72",x"72",x"6F",x"72",x"20",x"00",x"8D",x"1C",x"34",x"40",x"DE",x"3E",x"33",x"41",x"9E",
    x"40",x"30",x"01",x"A6",x"82",x"A7",x"C2",x"9C",x"44",x"26",x"F8",x"DF",x"42",x"35",x"C0",x"4F",
    x"58",x"D3",x"17",x"25",x"17",x"C3",x"00",x"3A",x"25",x"12",x"10",x"DF",x"11",x"10",x"93",x"11",
    x"22",x"0A",x"39",x"8E",x"C2",x"D2",x"BD",x"CD",x"E8",x"7E",x"CE",x"2C",x"C6",x"07",x"9E",x"19",
    x"30",x"1F",x"9F",x"72",x"D7",x"6F",x"86",x"11",x"97",x"79",x"BD",x"E1",x"96",x"0F",x"79",x"BD",
    x"EC",x"1E",x"DE",x"24",x"DF",x"70",x"9E",x"A7",x"27",x"04",x"96",x"A9",x"A7",x"84",x"BD",x"22",
    x"81",x"96",x"9E",x"27",x"03",x"BD",x"C4",x"24",x"10",x"DE",x"72",x"BD",x"C4",x"80",x"9E",x"2C",
    x"9F",x"74",x"DE",x"70",x"31",x"41",x"27",x"0E",x"DF",x"26",x"9F",x"2A",x"9E",x"21",x"27",x"06",
    x"96",x"23",x"10",x"27",x"1B",x"D4",x"8E",x"C2",x"DF",x"8D",x"AB",x"86",x"07",x"9D",x"E3",x"D6",
    x"6F",x"4F",x"BD",x"D8",x"3E",x"96",x"24",x"4C",x"27",x"03",x"BD",x"D8",x"37",x"0F",x"79",x"8D",
    x"92",x"BD",x"22",x"78",x"BD",x"EC",x"CF",x"25",x"F8",x"0D",x"7A",x"10",x"26",x"1F",x"73",x"9F",
    x"B3",x"9D",x"AC",x"27",x"EC",x"8E",x"FF",x"FF",x"9F",x"24",x"25",x"0E",x"C6",x"38",x"96",x"79",
    x"26",x"82",x"9E",x"B3",x"BD",x"DE",x"3A",x"7E",x"DF",x"5A",x"BD",x"C6",x"4B",x"BD",x"E1",x"07",
    x"9E",x"28",x"BF",x"24",x"4F",x"7F",x"24",x"51",x"9E",x"B3",x"A6",x"82",x"81",x"20",x"27",x"FA",
    x"30",x"01",x"A6",x"84",x"81",x"20",x"26",x"02",x"30",x"01",x"BD",x"DE",x"3A",x"34",x"06",x"8D",
    x"40",x"25",x"03",x"BD",x"CE",x"D9",x"B6",x"24",x"51",x"27",x"1A",x"DC",x"15",x"DD",x"40",x"E3",
    x"E1",x"DD",x"3E",x"BD",x"C2",x"E7",x"CE",x"24",x"4D",x"A6",x"C0",x"A7",x"80",x"9C",x"42",x"26",
    x"F8",x"9E",x"3E",x"9F",x"15",x"8D",x"02",x"20",x"88",x"8D",x"39",x"9E",x"44",x"EC",x"84",x"27",
    x"0F",x"33",x"04",x"A6",x"C0",x"26",x"FC",x"EF",x"84",x"AE",x"84",x"20",x"F0",x"43",x"9F",x"44",
    x"39",x"DC",x"28",x"9E",x"13",x"EE",x"84",x"27",x"F4",x"10",x"A3",x"02",x"23",x"F0",x"AE",x"84",
    x"20",x"F3",x"26",x"EA",x"0F",x"7F",x"9E",x"13",x"33",x"02",x"5F",x"6F",x"80",x"5A",x"26",x"FB",
    x"DF",x"15",x"0F",x"6E",x"9E",x"13",x"BD",x"C5",x"BD",x"BD",x"22",x"8D",x"BD",x"EA",x"08",x"8E",
    x"24",x"2B",x"CC",x"04",x"1A",x"A7",x"80",x"5A",x"26",x"FB",x"4F",x"97",x"23",x"DD",x"21",x"FD",
    x"25",x"81",x"FD",x"25",x"83",x"9E",x"1F",x"9F",x"1B",x"30",x"01",x"BF",x"20",x"70",x"8D",x"37",
    x"9E",x"15",x"9F",x"17",x"8E",x"80",x"4F",x"BF",x"24",x"27",x"8E",x"C7",x"52",x"BF",x"24",x"29",
    x"35",x"16",x"10",x"DE",x"19",x"6F",x"E2",x"10",x"DF",x"72",x"0F",x"2A",x"0F",x"2B",x"34",x"16",
    x"8E",x"25",x"85",x"9F",x"06",x"0F",x"9E",x"7E",x"CB",x"BD",x"27",x"0B",x"BD",x"C6",x"4B",x"BD",
    x"C4",x"11",x"24",x"05",x"7E",x"C5",x"D6",x"9E",x"13",x"30",x"1F",x"9F",x"30",x"39",x"BD",x"E1",
    x"C6",x"9D",x"B2",x"20",x"04",x"0F",x"79",x"1A",x"01",x"26",x"32",x"9E",x"B3",x"9F",x"2C",x"10",
    x"DE",x"72",x"06",x"A6",x"DE",x"24",x"30",x"41",x"27",x"06",x"DF",x"26",x"9E",x"2C",x"9F",x"2A",
    x"8E",x"C2",x"D7",x"0D",x"A6",x"10",x"2A",x"FE",x"B4",x"BD",x"CE",x"2C",x"7E",x"C3",x"75",x"C6",
    x"11",x"9E",x"2A",x"26",x"02",x"0E",x"FB",x"9F",x"B3",x"9E",x"26",x"9F",x"24",x"39",x"27",x"5E",
    x"DC",x"1F",x"93",x"19",x"34",x"0E",x"9D",x"B2",x"81",x"2C",x"27",x"05",x"BD",x"C9",x"85",x"ED",
    x"E4",x"BD",x"EA",x"22",x"34",x"10",x"9D",x"B2",x"27",x"11",x"9D",x"C2",x"81",x"2C",x"27",x"0B",
    x"BD",x"CC",x"BA",x"30",x"1F",x"9C",x"A1",x"22",x"3F",x"AF",x"E4",x"D6",x"AA",x"9D",x"B2",x"27",
    x"09",x"BD",x"CC",x"AB",x"C1",x"80",x"10",x"22",x"5C",x"DC",x"E7",x"64",x"86",x"08",x"3D",x"DD",
    x"4E",x"35",x"06",x"93",x"4E",x"1F",x"01",x"A3",x"E1",x"25",x"1D",x"1F",x"03",x"83",x"00",x"3A",
    x"25",x"16",x"93",x"15",x"25",x"12",x"DF",x"19",x"9F",x"1F",x"35",x"04",x"D7",x"AA",x"35",x"10",
    x"10",x"DE",x"19",x"34",x"10",x"7E",x"C4",x"39",x"7E",x"C3",x"1C",x"81",x"22",x"10",x"27",x"1D",
    x"02",x"BD",x"E1",x"C6",x"9D",x"B2",x"10",x"27",x"FE",x"DA",x"BD",x"C4",x"39",x"20",x"19",x"1F",
    x"89",x"9D",x"AC",x"C1",x"BB",x"27",x"3F",x"C1",x"BC",x"26",x"6F",x"C6",x"03",x"BD",x"C2",x"FF",
    x"DE",x"B3",x"9E",x"24",x"86",x"BC",x"34",x"52",x"8D",x"2C",x"7E",x"DF",x"26",x"C6",x"3A",x"21",
    x"5F",x"9E",x"B3",x"0F",x"00",x"1E",x"89",x"D6",x"00",x"97",x"00",x"A6",x"84",x"27",x"5A",x"91",
    x"00",x"27",x"56",x"30",x"01",x"81",x"22",x"27",x"EC",x"4C",x"26",x"02",x"30",x"01",x"81",x"8A",
    x"26",x"E9",x"0C",x"62",x"20",x"E5",x"9D",x"B2",x"BD",x"C6",x"4B",x"8D",x"D3",x"30",x"01",x"DC",
    x"28",x"10",x"93",x"24",x"22",x"02",x"9E",x"13",x"BD",x"C4",x"15",x"25",x"19",x"30",x"1F",x"20",
    x"26",x"26",x"26",x"86",x"FF",x"97",x"3B",x"BD",x"CF",x"63",x"32",x"84",x"10",x"DF",x"72",x"81",
    x"3B",x"27",x"09",x"C6",x"03",x"8C",x"C6",x"08",x"0E",x"FB",x"0E",x"F9",x"35",x"52",x"9F",x"24",
    x"DF",x"B3",x"8D",x"99",x"8C",x"8D",x"99",x"9F",x"B3",x"39",x"9D",x"D9",x"9D",x"B2",x"81",x"87",
    x"26",x"0A",x"9D",x"AC",x"9D",x"CA",x"81",x"BB",x"27",x"06",x"0E",x"F9",x"C6",x"C4",x"9D",x"E0",
    x"BD",x"D5",x"83",x"26",x"13",x"0F",x"62",x"8D",x"D9",x"4D",x"27",x"DD",x"9D",x"AC",x"81",x"8F",
    x"26",x"F5",x"0A",x"62",x"2A",x"F1",x"9D",x"AC",x"9D",x"B2",x"25",x"8C",x"7E",x"DF",x"60",x"81",
    x"98",x"27",x"66",x"BD",x"22",x"72",x"9D",x"E6",x"C6",x"87",x"9D",x"E0",x"34",x"02",x"81",x"BC",
    x"27",x"04",x"81",x"BB",x"26",x"C4",x"0A",x"4F",x"26",x"05",x"35",x"04",x"7E",x"C5",x"61",x"9D",
    x"AC",x"8D",x"08",x"81",x"2C",x"27",x"EF",x"9D",x"B2",x"35",x"84",x"9E",x"FE",x"9F",x"28",x"25",
    x"02",x"0E",x"B2",x"80",x"30",x"97",x"00",x"DC",x"28",x"81",x"18",x"22",x"9D",x"58",x"49",x"58",
    x"49",x"D3",x"28",x"58",x"49",x"DB",x"00",x"89",x"00",x"DD",x"28",x"9D",x"AC",x"20",x"E0",x"9D",
    x"F0",x"9F",x"3B",x"BD",x"CF",x"88",x"9D",x"C5",x"10",x"26",x"11",x"75",x"BD",x"CB",x"F9",x"BD",
    x"EF",x"EF",x"DE",x"3B",x"E7",x"C4",x"AF",x"41",x"39",x"9D",x"AC",x"C6",x"87",x"9D",x"E0",x"C6",
    x"BB",x"9D",x"E0",x"8D",x"B6",x"9E",x"28",x"27",x"0A",x"BD",x"C4",x"11",x"10",x"25",x"FF",x"36",
    x"9F",x"21",x"39",x"9F",x"21",x"96",x"23",x"27",x"F9",x"9E",x"70",x"9F",x"24",x"7E",x"C3",x"48",
    x"6E",x"9F",x"22",x"13",x"9D",x"AC",x"1F",x"89",x"58",x"9D",x"AC",x"C1",x"4C",x"22",x"F1",x"34",
    x"04",x"C1",x"3E",x"24",x"0A",x"8D",x"68",x"E6",x"E4",x"C1",x"34",x"24",x"02",x"8D",x"5C",x"35",
    x"04",x"BE",x"22",x"09",x"6E",x"95",x"4F",x"D6",x"6F",x"8C",x"DC",x"70",x"BD",x"D8",x"45",x"0E",
    x"AC",x"9E",x"B3",x"BD",x"CB",x"6F",x"9E",x"5E",x"9F",x"B3",x"39",x"9D",x"AC",x"27",x"4F",x"24",
    x"05",x"9D",x"CA",x"7E",x"D1",x"E3",x"BD",x"C8",x"A1",x"24",x"12",x"9D",x"F0",x"9F",x"4E",x"9D",
    x"C5",x"27",x"E7",x"7E",x"D6",x"8D",x"86",x"7D",x"8D",x"39",x"7E",x"D2",x"8F",x"8E",x"C0",x"4E",
    x"A1",x"81",x"22",x"FC",x"10",x"26",x"5B",x"21",x"E6",x"1F",x"8E",x"C7",x"06",x"6E",x"85",x"86",
    x"5A",x"8D",x"20",x"BD",x"D6",x"27",x"7E",x"C8",x"69",x"8D",x"04",x"9D",x"D9",x"0E",x"DE",x"C6",
    x"28",x"8C",x"C6",x"2C",x"E1",x"9F",x"21",x"B3",x"26",x"02",x"0E",x"AC",x"0E",x"F9",x"C6",x"16",
    x"0E",x"FB",x"4F",x"34",x"02",x"C6",x"01",x"BD",x"C2",x"FF",x"8D",x"9F",x"9D",x"B2",x"80",x"C7",
    x"25",x"10",x"81",x"0E",x"22",x"0C",x"C6",x"03",x"3D",x"8E",x"C0",x"67",x"A6",x"85",x"A1",x"E4",
    x"22",x"02",x"35",x"82",x"97",x"3D",x"5C",x"EE",x"85",x"C6",x"04",x"D7",x"42",x"EC",x"9F",x"21",
    x"B3",x"8E",x"C0",x"92",x"30",x"02",x"0A",x"42",x"27",x"09",x"10",x"A3",x"81",x"26",x"F5",x"EE",
    x"84",x"9D",x"AC",x"34",x"40",x"8D",x"5C",x"96",x"3D",x"8D",x"B8",x"97",x"3D",x"8D",x"60",x"96",
    x"3D",x"D6",x"57",x"C1",x"03",x"27",x"2F",x"4C",x"2B",x"14",x"81",x"51",x"23",x"1E",x"80",x"7B",
    x"44",x"27",x"19",x"96",x"4B",x"44",x"25",x"24",x"9B",x"57",x"81",x"04",x"25",x"06",x"9D",x"E9",
    x"8D",x"55",x"9D",x"E9",x"8D",x"51",x"35",x"10",x"AD",x"84",x"20",x"90",x"BD",x"D6",x"27",x"8D",
    x"46",x"BD",x"D6",x"27",x"20",x"F0",x"97",x"3D",x"9D",x"C5",x"27",x"03",x"7E",x"D6",x"5C",x"8D",
    x"36",x"86",x"64",x"91",x"3D",x"27",x"DF",x"8E",x"D2",x"AC",x"AC",x"E1",x"26",x"EE",x"8E",x"CB",
    x"C2",x"20",x"D5",x"35",x"20",x"DC",x"4B",x"9E",x"4D",x"DE",x"4F",x"34",x"56",x"6E",x"A4",x"35",
    x"20",x"35",x"56",x"DF",x"5B",x"9F",x"59",x"DD",x"57",x"6E",x"A4",x"35",x"20",x"35",x"56",x"DF",
    x"4F",x"9F",x"4D",x"DD",x"4B",x"6E",x"A4",x"DC",x"58",x"9E",x"4C",x"9F",x"58",x"DD",x"4C",x"96",
    x"5C",x"D6",x"50",x"D7",x"5C",x"97",x"50",x"96",x"4B",x"D6",x"57",x"97",x"57",x"D7",x"4B",x"9E",
    x"4E",x"BD",x"D6",x"7B",x"9F",x"5A",x"39",x"BD",x"CB",x"FC",x"BD",x"CB",x"F0",x"BD",x"CB",x"F9",
    x"D1",x"53",x"27",x"06",x"4A",x"25",x"03",x"D6",x"53",x"40",x"97",x"50",x"DE",x"54",x"5C",x"5A",
    x"27",x"0C",x"A6",x"80",x"A1",x"C0",x"27",x"F7",x"C6",x"01",x"24",x"04",x"50",x"8C",x"D6",x"50",
    x"1D",x"20",x"0B",x"9D",x"C5",x"27",x"D0",x"2A",x"02",x"8D",x"C4",x"BD",x"D5",x"B7",x"DD",x"4E",
    x"4F",x"5F",x"9E",x"4E",x"39",x"8D",x"EC",x"26",x"02",x"43",x"53",x"0E",x"ED",x"8D",x"E4",x"2B",
    x"F8",x"20",x"F8",x"8D",x"DE",x"27",x"F2",x"20",x"F6",x"8D",x"F2",x"8C",x"8D",x"E7",x"8C",x"8D",
    x"F2",x"03",x"4E",x"03",x"4F",x"39",x"94",x"5A",x"D4",x"5B",x"20",x"DF",x"9A",x"5A",x"DA",x"5B",
    x"20",x"D9",x"98",x"5A",x"D8",x"5B",x"20",x"D3",x"43",x"53",x"20",x"F0",x"12",x"8D",x"F3",x"20",
    x"C8",x"81",x"5B",x"24",x"04",x"80",x"41",x"80",x"BF",x"39",x"0F",x"3A",x"DE",x"B3",x"DF",x"34",
    x"A6",x"C0",x"8D",x"ED",x"25",x"02",x"0E",x"F9",x"5F",x"A6",x"C0",x"C1",x"0F",x"27",x"01",x"5C",
    x"8D",x"DF",x"25",x"F5",x"9D",x"B9",x"25",x"F1",x"D7",x"36",x"DF",x"B3",x"8E",x"C0",x"62",x"80",
    x"21",x"81",x"04",x"23",x"09",x"9D",x"CA",x"8E",x"23",x"EA",x"A6",x"9F",x"21",x"34",x"E6",x"86",
    x"27",x"F3",x"0D",x"3A",x"2B",x"0A",x"26",x"06",x"9D",x"B2",x"81",x"28",x"26",x"02",x"CB",x"08",
    x"D7",x"4B",x"9E",x"15",x"9C",x"17",x"27",x"57",x"8D",x"43",x"E6",x"84",x"54",x"54",x"54",x"54",
    x"D7",x"39",x"E6",x"84",x"C4",x"0F",x"A1",x"80",x"27",x"14",x"3A",x"4F",x"8D",x"3C",x"27",x"02",
    x"EC",x"81",x"30",x"8B",x"20",x"DE",x"96",x"3A",x"84",x"80",x"AA",x"C0",x"5A",x"39",x"8D",x"F6",
    x"2A",x"E4",x"8D",x"26",x"27",x"3A",x"96",x"3A",x"26",x"64",x"8D",x"7B",x"A1",x"80",x"26",x"64",
    x"EC",x"E1",x"BD",x"C9",x"E1",x"0A",x"02",x"26",x"F7",x"30",x"8B",x"20",x"23",x"DE",x"34",x"96",
    x"4B",x"48",x"48",x"48",x"48",x"9B",x"36",x"D6",x"36",x"39",x"D6",x"39",x"C5",x"08",x"39",x"D6",
    x"4B",x"D7",x"39",x"0D",x"3A",x"2E",x"0B",x"8D",x"F1",x"26",x"3D",x"8D",x"0E",x"10",x"9F",x"17",
    x"9F",x"37",x"39",x"86",x"01",x"97",x"3A",x"BD",x"C8",x"AC",x"5F",x"9E",x"17",x"4F",x"DB",x"36",
    x"5C",x"31",x"8B",x"BD",x"C3",x"05",x"8D",x"C5",x"A7",x"80",x"8D",x"9A",x"2A",x"FA",x"6F",x"84",
    x"6F",x"01",x"39",x"9D",x"AC",x"9D",x"CD",x"BD",x"D6",x"27",x"2A",x"F6",x"0E",x"F6",x"44",x"26",
    x"F1",x"C6",x"0A",x"8C",x"C6",x"09",x"0E",x"FB",x"DE",x"34",x"34",x"40",x"8D",x"CC",x"BD",x"CA",
    x"25",x"35",x"40",x"DF",x"B3",x"0E",x"F0",x"35",x"20",x"D6",x"39",x"C4",x"07",x"4F",x"DE",x"3A",
    x"34",x"76",x"8D",x"CF",x"35",x"76",x"DF",x"3A",x"4C",x"2B",x"D1",x"DE",x"4E",x"34",x"42",x"97",
    x"02",x"9D",x"B2",x"81",x"2C",x"35",x"02",x"27",x"E5",x"D7",x"39",x"9D",x"DE",x"33",x"84",x"30",
    x"02",x"4F",x"5F",x"DD",x"5E",x"5C",x"DD",x"60",x"96",x"02",x"6E",x"A4",x"ED",x"84",x"83",x"00",
    x"01",x"8D",x"2A",x"D3",x"5E",x"2B",x"AD",x"DD",x"5E",x"EC",x"81",x"8D",x"25",x"DD",x"60",x"DC",
    x"5E",x"DD",x"4E",x"D6",x"39",x"96",x"4E",x"3D",x"D7",x"4E",x"2B",x"98",x"4D",x"26",x"95",x"96",
    x"4F",x"D6",x"39",x"D7",x"4B",x"3D",x"9B",x"4E",x"2B",x"8A",x"DD",x"4E",x"39",x"10",x"A3",x"84",
    x"24",x"82",x"DD",x"5A",x"DC",x"60",x"9D",x"ED",x"BD",x"D2",x"F2",x"9D",x"C5",x"2A",x"DE",x"DC",
    x"4E",x"39",x"BD",x"C9",x"63",x"8D",x"80",x"A7",x"80",x"1F",x"89",x"48",x"4C",x"A7",x"41",x"6F",
    x"C4",x"BD",x"C2",x"FF",x"EC",x"E1",x"C3",x"00",x"01",x"0D",x"3A",x"26",x"03",x"CC",x"00",x"0B",
    x"8D",x"9A",x"0A",x"02",x"26",x"EE",x"DB",x"4B",x"89",x"00",x"DD",x"4E",x"E3",x"C4",x"ED",x"C1",
    x"BD",x"C3",x"01",x"10",x"9E",x"4E",x"6F",x"80",x"31",x"3F",x"26",x"FA",x"9F",x"17",x"39",x"9D",
    x"AC",x"8D",x"BF",x"9D",x"B2",x"81",x"2C",x"27",x"F6",x"39",x"9D",x"C5",x"26",x"0B",x"BD",x"CB",
    x"F9",x"8D",x"4B",x"DC",x"1B",x"93",x"19",x"20",x"04",x"1F",x"40",x"93",x"17",x"7E",x"D8",x"45",
    x"0F",x"03",x"4F",x"34",x"06",x"DC",x"1B",x"A3",x"E0",x"1F",x"01",x"9C",x"19",x"25",x"23",x"9F",
    x"1B",x"30",x"01",x"9F",x"1D",x"35",x"84",x"6D",x"1F",x"2B",x"14",x"A6",x"84",x"27",x"10",x"EC",
    x"01",x"10",x"93",x"1B",x"22",x"09",x"10",x"93",x"44",x"23",x"04",x"9F",x"46",x"DD",x"44",x"30",
    x"03",x"39",x"C6",x"0E",x"03",x"03",x"27",x"78",x"8D",x"04",x"35",x"04",x"20",x"C4",x"9E",x"1F",
    x"9F",x"1B",x"4F",x"5F",x"DD",x"46",x"9E",x"19",x"9F",x"44",x"8E",x"25",x"85",x"9C",x"06",x"27",
    x"04",x"8D",x"C8",x"20",x"F8",x"4F",x"9E",x"15",x"30",x"86",x"9C",x"17",x"27",x"33",x"E6",x"80",
    x"1F",x"98",x"C4",x"0F",x"3A",x"44",x"44",x"44",x"44",x"85",x"08",x"26",x"08",x"81",x"03",x"26",
    x"E7",x"8D",x"A4",x"20",x"E5",x"81",x"0B",x"27",x"06",x"EC",x"81",x"30",x"8B",x"20",x"DB",x"EC",
    x"81",x"33",x"8B",x"DF",x"3E",x"E6",x"80",x"58",x"3A",x"9C",x"3E",x"27",x"CD",x"8D",x"8C",x"20",
    x"F8",x"9E",x"46",x"27",x"9C",x"4F",x"E6",x"84",x"5A",x"D3",x"44",x"DD",x"40",x"9E",x"1B",x"9F",
    x"3E",x"BD",x"C2",x"E9",x"DE",x"46",x"9E",x"42",x"AF",x"41",x"30",x"1F",x"20",x"92",x"C6",x"10",
    x"0E",x"FB",x"4F",x"5F",x"DD",x"00",x"9F",x"60",x"9F",x"54",x"C6",x"FF",x"5C",x"A6",x"80",x"27",
    x"0C",x"91",x"00",x"27",x"04",x"91",x"01",x"26",x"F3",x"81",x"22",x"27",x"02",x"30",x"1F",x"9F",
    x"5E",x"96",x"01",x"81",x"2C",x"26",x"0A",x"5C",x"5A",x"27",x"06",x"A6",x"82",x"81",x"20",x"27",
    x"F7",x"D7",x"53",x"39",x"9D",x"D1",x"BD",x"D8",x"52",x"8D",x"C7",x"20",x"12",x"30",x"1F",x"86",
    x"22",x"1F",x"89",x"30",x"01",x"8D",x"BD",x"DE",x"60",x"11",x"83",x"25",x"54",x"22",x"06",x"8D",
    x"6C",x"9E",x"60",x"8D",x"4B",x"9E",x"06",x"8C",x"25",x"A3",x"27",x"A2",x"86",x"03",x"97",x"4B",
    x"9F",x"08",x"9F",x"4E",x"96",x"53",x"A7",x"80",x"DE",x"54",x"EF",x"81",x"9F",x"06",x"39",x"8D",
    x"56",x"10",x"27",x"0A",x"36",x"DE",x"B3",x"9F",x"B3",x"3A",x"A6",x"84",x"97",x"A9",x"9F",x"A7",
    x"34",x"52",x"6F",x"84",x"BD",x"C6",x"F1",x"35",x"52",x"A7",x"84",x"DF",x"B3",x"4F",x"5F",x"DD",
    x"A7",x"39",x"E6",x"9F",x"21",x"5A",x"9E",x"4E",x"EB",x"84",x"24",x"13",x"C6",x"0F",x"0E",x"FB",
    x"DE",x"1D",x"5C",x"20",x"04",x"A6",x"80",x"A7",x"C0",x"5A",x"26",x"F9",x"DF",x"1D",x"39",x"8D",
    x"0C",x"8D",x"19",x"8D",x"14",x"8D",x"E9",x"8D",x"13",x"8D",x"E5",x"20",x"98",x"BD",x"CA",x"80",
    x"9F",x"54",x"D7",x"53",x"39",x"9D",x"D9",x"9D",x"D6",x"DE",x"4E",x"8C",x"DE",x"5A",x"11",x"93",
    x"08",x"26",x"06",x"DF",x"06",x"30",x"5D",x"9F",x"08",x"AE",x"41",x"E6",x"C4",x"39",x"8D",x"07",
    x"8C",x"8D",x"E4",x"0E",x"EC",x"9D",x"D9",x"8D",x"DE",x"27",x"73",x"E6",x"84",x"39",x"8D",x"70",
    x"96",x"80",x"90",x"4F",x"8C",x"8D",x"69",x"D1",x"80",x"23",x"03",x"4F",x"D6",x"80",x"34",x"06",
    x"9C",x"13",x"25",x"04",x"9C",x"15",x"25",x"02",x"8D",x"B3",x"DE",x"82",x"8D",x"C0",x"35",x"04",
    x"3A",x"35",x"04",x"9C",x"13",x"25",x"04",x"9C",x"15",x"25",x"03",x"7E",x"CB",x"83",x"8D",x"A0",
    x"20",x"99",x"8D",x"5E",x"CB",x"80",x"25",x"36",x"D7",x"4F",x"8C",x"8D",x"55",x"C6",x"01",x"8D",
    x"8C",x"96",x"4F",x"A7",x"84",x"20",x"E9",x"8D",x"2E",x"D7",x"81",x"27",x"21",x"C6",x"FF",x"D7",
    x"4F",x"9D",x"B2",x"81",x"29",x"27",x"02",x"8D",x"32",x"9D",x"DE",x"0A",x"81",x"96",x"81",x"D6",
    x"80",x"D0",x"81",x"24",x"01",x"5F",x"D1",x"4F",x"23",x"A4",x"D6",x"4F",x"20",x"A0",x"0E",x"F6",
    x"8D",x"05",x"9D",x"DE",x"DC",x"4E",x"39",x"8D",x"0A",x"DE",x"4E",x"34",x"40",x"8D",x"0C",x"7E",
    x"FF",x"DB",x"12",x"9D",x"D9",x"0E",x"D6",x"8D",x"11",x"9F",x"28",x"9D",x"C2",x"8C",x"9D",x"AC",
    x"9D",x"CD",x"BD",x"C9",x"87",x"4D",x"26",x"D6",x"0E",x"B2",x"9D",x"CD",x"9D",x"E9",x"96",x"50",
    x"2A",x"06",x"8E",x"CD",x"46",x"BD",x"D3",x"99",x"96",x"4C",x"81",x"90",x"22",x"C0",x"BD",x"D5",
    x"EE",x"9E",x"4E",x"39",x"BD",x"E1",x"01",x"8D",x"E3",x"E6",x"84",x"0E",x"EC",x"BD",x"E1",x"01",
    x"8D",x"C5",x"9E",x"28",x"E7",x"84",x"39",x"9D",x"D9",x"C6",x"01",x"34",x"04",x"9D",x"C5",x"27",
    x"0A",x"8D",x"BF",x"E7",x"E4",x"27",x"97",x"9D",x"C2",x"8D",x"A8",x"DC",x"4E",x"34",x"06",x"9D",
    x"C2",x"BD",x"C7",x"2B",x"BD",x"CB",x"F7",x"9F",x"5E",x"D7",x"64",x"35",x"40",x"BD",x"CB",x"FE",
    x"D7",x"63",x"35",x"04",x"D7",x"62",x"D1",x"63",x"22",x"29",x"0D",x"64",x"27",x"22",x"5A",x"3A",
    x"9F",x"60",x"DE",x"5E",x"96",x"63",x"90",x"62",x"4C",x"91",x"64",x"25",x"16",x"D6",x"64",x"A6",
    x"80",x"A1",x"C0",x"27",x"08",x"0C",x"62",x"9E",x"60",x"30",x"01",x"20",x"E3",x"5A",x"26",x"EF",
    x"D6",x"62",x"21",x"5F",x"0E",x"EC",x"91",x"00",x"00",x"00",x"9D",x"DB",x"BD",x"D6",x"27",x"9D",
    x"DE",x"9D",x"CA",x"4F",x"5F",x"0D",x"4E",x"2A",x"02",x"DD",x"4E",x"4C",x"DD",x"5A",x"9D",x"F3",
    x"27",x"06",x"0F",x"5A",x"96",x"7E",x"97",x"5B",x"4F",x"BD",x"D3",x"77",x"D6",x"4F",x"D0",x"7D",
    x"24",x"05",x"BD",x"CD",x"F0",x"D6",x"4F",x"7E",x"CE",x"19",x"27",x"74",x"8D",x"03",x"0F",x"79",
    x"39",x"81",x"23",x"26",x"0C",x"BD",x"E1",x"D0",x"BD",x"E4",x"16",x"9D",x"B2",x"27",x"61",x"9D",
    x"C2",x"81",x"BF",x"10",x"27",x"03",x"4B",x"26",x"01",x"39",x"81",x"BA",x"27",x"AC",x"81",x"BE",
    x"27",x"70",x"81",x"2C",x"27",x"55",x"81",x"3B",x"27",x"77",x"9D",x"D9",x"9D",x"C5",x"34",x"02",
    x"27",x"06",x"BD",x"D8",x"52",x"BD",x"CB",x"6D",x"9D",x"F3",x"DC",x"7D",x"3D",x"27",x"0A",x"9E",
    x"4E",x"AB",x"84",x"91",x"7E",x"23",x"02",x"8D",x"27",x"8D",x"64",x"35",x"02",x"0D",x"8F",x"27",
    x"06",x"8D",x"71",x"9D",x"B2",x"20",x"C0",x"4D",x"27",x"08",x"9D",x"B2",x"81",x"2C",x"27",x"02",
    x"8D",x"5C",x"9D",x"B2",x"26",x"B4",x"20",x"08",x"9D",x"F3",x"27",x"04",x"96",x"7D",x"27",x"A9",
    x"8D",x"52",x"86",x"0A",x"9D",x"F3",x"0D",x"8F",x"27",x"4C",x"39",x"9D",x"F3",x"27",x"0A",x"D6",
    x"7D",x"D1",x"7C",x"25",x"06",x"D0",x"7E",x"20",x"06",x"D6",x"7D",x"D0",x"7B",x"24",x"FC",x"50",
    x"20",x"07",x"BD",x"CC",x"AE",x"81",x"29",x"26",x"2F",x"9D",x"F3",x"0D",x"8F",x"26",x"02",x"8D",
    x"07",x"9D",x"AC",x"20",x"B0",x"8D",x"17",x"5A",x"5D",x"26",x"FA",x"39",x"BD",x"CB",x"6F",x"BD",
    x"CB",x"F9",x"5C",x"5A",x"27",x"B8",x"A6",x"80",x"8D",x"0C",x"20",x"F7",x"8D",x"03",x"86",x"20",
    x"8C",x"86",x"3F",x"8C",x"86",x"0D",x"0E",x"E3",x"0E",x"F9",x"96",x"79",x"26",x"07",x"C6",x"18",
    x"3F",x"02",x"BD",x"E4",x"79",x"BD",x"CD",x"F0",x"9C",x"69",x"26",x"06",x"BD",x"E1",x"96",x"7E",
    x"C3",x"7D",x"9F",x"67",x"EC",x"02",x"BD",x"D8",x"3E",x"BD",x"CE",x"3E",x"9E",x"67",x"BD",x"DD",
    x"DA",x"8E",x"24",x"52",x"A6",x"80",x"27",x"04",x"9D",x"E3",x"20",x"F8",x"9E",x"67",x"AE",x"84",
    x"20",x"C8",x"4F",x"5F",x"DD",x"67",x"8E",x"F9",x"FF",x"9F",x"69",x"9D",x"B2",x"27",x"1C",x"8D",
    x"2F",x"9E",x"28",x"9F",x"67",x"9D",x"B2",x"26",x"04",x"9F",x"69",x"20",x"0E",x"C6",x"C8",x"9D",
    x"E0",x"27",x"08",x"8D",x"1B",x"8D",x"2C",x"9E",x"28",x"9F",x"69",x"9E",x"69",x"9C",x"67",x"25",
    x"16",x"30",x"01",x"9F",x"28",x"8D",x"06",x"9F",x"69",x"9E",x"67",x"9F",x"28",x"7E",x"C4",x"11",
    x"9D",x"B2",x"7E",x"C6",x"4B",x"26",x"02",x"0E",x"F6",x"8D",x"B7",x"8D",x"0A",x"BD",x"C3",x"F9",
    x"7E",x"C3",x"7D",x"27",x"13",x"0E",x"F9",x"DE",x"69",x"9F",x"44",x"11",x"93",x"15",x"27",x"06",
    x"A6",x"C0",x"A7",x"80",x"20",x"F5",x"9F",x"15",x"39",x"C6",x"04",x"8C",x"C6",x"03",x"8C",x"C6",
    x"02",x"D7",x"3D",x"8D",x"21",x"8E",x"23",x"EA",x"3A",x"34",x"04",x"81",x"C8",x"26",x"02",x"8D",
    x"13",x"E0",x"E0",x"2B",x"D0",x"96",x"3D",x"A7",x"80",x"5A",x"2A",x"FB",x"9D",x"B2",x"27",x"D8",
    x"9D",x"C2",x"20",x"DF",x"9D",x"AC",x"BD",x"C8",x"A1",x"24",x"BA",x"1F",x"89",x"0E",x"AC",x"86",
    x"4F",x"97",x"6E",x"39",x"9D",x"E6",x"26",x"FB",x"5D",x"27",x"9C",x"0E",x"FB",x"C6",x"14",x"0D",
    x"23",x"27",x"F8",x"0F",x"6F",x"81",x"82",x"27",x"1B",x"9D",x"B2",x"24",x"0A",x"BD",x"C6",x"4B",
    x"26",x"11",x"BD",x"C5",x"AB",x"20",x"0A",x"8D",x"8A",x"9E",x"70",x"9F",x"24",x"9E",x"74",x"9F",
    x"B3",x"0F",x"23",x"39",x"9D",x"AC",x"8D",x"EF",x"6D",x"80",x"26",x"02",x"30",x"03",x"9F",x"B3",
    x"7E",x"C5",x"E2",x"30",x"64",x"9F",x"0A",x"A6",x"84",x"C6",x"13",x"80",x"81",x"26",x"15",x"AE",
    x"01",x"9F",x"0C",x"9E",x"3B",x"27",x"09",x"9C",x"0C",x"27",x"09",x"9E",x"0A",x"3A",x"20",x"E5",
    x"9E",x"0C",x"9F",x"3B",x"9E",x"0A",x"4D",x"39",x"C6",x"D4",x"9D",x"E0",x"96",x"4B",x"34",x"02",
    x"9D",x"D9",x"35",x"02",x"7E",x"D6",x"65",x"9D",x"F0",x"9F",x"3B",x"9D",x"D1",x"8D",x"E9",x"8E",
    x"21",x"65",x"BD",x"D7",x"F3",x"32",x"62",x"BD",x"C5",x"7D",x"9F",x"6C",x"1F",x"41",x"BD",x"CF",
    x"65",x"3A",x"26",x"0A",x"EC",x"1E",x"93",x"6C",x"26",x"F4",x"32",x"84",x"9F",x"72",x"C6",x"0A",
    x"BD",x"C2",x"FF",x"9E",x"6C",x"DC",x"24",x"34",x"16",x"C6",x"BB",x"8D",x"BD",x"32",x"7C",x"1F",
    x"41",x"BD",x"D7",x"F7",x"8E",x"00",x"01",x"9F",x"4E",x"9D",x"C5",x"2B",x"06",x"8E",x"DC",x"33",
    x"BD",x"D6",x"8D",x"9D",x"B2",x"81",x"C6",x"26",x"04",x"9D",x"AC",x"8D",x"9F",x"BD",x"D5",x"83",
    x"D7",x"50",x"BD",x"C7",x"E3",x"9D",x"B2",x"BD",x"CE",x"D3",x"5F",x"9E",x"24",x"9F",x"6C",x"9D",
    x"CA",x"5C",x"9D",x"AC",x"27",x"07",x"4C",x"26",x"1B",x"9D",x"AC",x"20",x"F5",x"4D",x"26",x"F2",
    x"9E",x"B3",x"EE",x"01",x"26",x"04",x"C6",x"17",x"0E",x"FB",x"30",x"03",x"EE",x"80",x"DF",x"6C",
    x"9F",x"B3",x"20",x"DE",x"81",x"82",x"27",x"D9",x"81",x"83",x"26",x"D6",x"5A",x"27",x"1C",x"9D",
    x"AC",x"27",x"DA",x"9E",x"6C",x"9F",x"24",x"34",x"04",x"9D",x"F0",x"35",x"04",x"AE",x"6A",x"9F",
    x"24",x"9D",x"B2",x"27",x"C8",x"81",x"2C",x"27",x"E3",x"0E",x"F9",x"9D",x"AC",x"DE",x"B3",x"9E",
    x"3B",x"86",x"81",x"34",x"52",x"9E",x"6C",x"9F",x"24",x"8D",x"00",x"86",x"4F",x"97",x"6B",x"9E",
    x"FE",x"9F",x"3B",x"9E",x"B3",x"9F",x"6C",x"9D",x"B2",x"27",x"04",x"9D",x"F0",x"9F",x"3B",x"BD",
    x"CF",x"63",x"27",x"04",x"C6",x"01",x"0E",x"FB",x"1F",x"14",x"AE",x"03",x"9C",x"6C",x"26",x"F4",
    x"A6",x"65",x"97",x"4B",x"97",x"57",x"96",x"6B",x"27",x"21",x"8E",x"21",x"65",x"BD",x"D6",x"8D",
    x"BD",x"D7",x"F1",x"30",x"6B",x"BD",x"D3",x"85",x"BD",x"D5",x"B7",x"EB",x"6A",x"27",x"27",x"AE",
    x"6F",x"9F",x"24",x"AE",x"E8",x"11",x"9F",x"B3",x"7E",x"DF",x"26",x"9E",x"3B",x"BD",x"D6",x"8D",
    x"30",x"66",x"BD",x"D3",x"85",x"E6",x"6A",x"D7",x"5C",x"96",x"4B",x"34",x"02",x"BD",x"D2",x"AC",
    x"96",x"4B",x"A1",x"E0",x"27",x"CA",x"32",x"E8",x"13",x"30",x"E4",x"9F",x"72",x"9D",x"B2",x"81",
    x"2C",x"26",x"D5",x"9D",x"AC",x"0F",x"6B",x"8D",x"88",x"9D",x"F0",x"9F",x"4E",x"BD",x"D6",x"51",
    x"0E",x"DE",x"9D",x"AC",x"BD",x"CB",x"F5",x"C6",x"3B",x"9D",x"E0",x"E6",x"C4",x"4F",x"34",x"14",
    x"97",x"78",x"5D",x"27",x"2B",x"0F",x"76",x"0F",x"77",x"A6",x"80",x"81",x"5E",x"27",x"1E",x"81",
    x"2B",x"26",x"04",x"86",x"08",x"20",x"06",x"81",x"2A",x"26",x"08",x"86",x"20",x"9A",x"78",x"97",
    x"78",x"20",x"0A",x"81",x"23",x"27",x"1F",x"81",x"2E",x"27",x"6F",x"9D",x"E3",x"5A",x"26",x"D9",
    x"35",x"14",x"9D",x"B2",x"10",x"27",x"FC",x"C8",x"81",x"3B",x"26",x"02",x"0E",x"AC",x"96",x"78",
    x"27",x"02",x"20",x"BA",x"0E",x"F6",x"0C",x"77",x"5A",x"27",x"12",x"A6",x"80",x"81",x"23",x"27",
    x"F5",x"81",x"2E",x"27",x"45",x"81",x"5E",x"26",x"02",x"0C",x"78",x"30",x"1F",x"96",x"78",x"85",
    x"08",x"27",x"02",x"0C",x"77",x"96",x"77",x"9B",x"76",x"81",x"18",x"24",x"D7",x"86",x"80",x"9A",
    x"78",x"97",x"78",x"9D",x"B2",x"27",x"B9",x"34",x"14",x"9D",x"CD",x"BD",x"D8",x"54",x"30",x"1F",
    x"BD",x"CE",x"2C",x"35",x"14",x"9D",x"B2",x"27",x"0C",x"81",x"3B",x"27",x"08",x"81",x"2C",x"10",
    x"26",x"50",x"76",x"9D",x"AC",x"86",x"80",x"16",x"FF",x"66",x"0C",x"76",x"5A",x"27",x"BE",x"A6",
    x"80",x"81",x"23",x"20",x"AE",x"9D",x"AC",x"9D",x"AC",x"81",x"48",x"26",x"45",x"9D",x"AC",x"25",
    x"0B",x"81",x"47",x"BD",x"C8",x"A3",x"10",x"24",x"06",x"9D",x"80",x"07",x"80",x"30",x"C6",x"04",
    x"08",x"4F",x"09",x"4E",x"10",x"25",x"03",x"26",x"5A",x"26",x"F5",x"9B",x"4F",x"97",x"4F",x"20",
    x"DC",x"81",x"02",x"26",x"08",x"96",x"4F",x"84",x"0F",x"27",x"02",x"9D",x"E9",x"BD",x"D4",x"B1",
    x"BD",x"D6",x"80",x"35",x"04",x"4F",x"BD",x"D2",x"C8",x"BD",x"D3",x"9B",x"20",x"15",x"96",x"4B",
    x"80",x"02",x"39",x"5F",x"BD",x"D5",x"DB",x"DD",x"44",x"DD",x"42",x"8D",x"4A",x"81",x"26",x"27",
    x"A4",x"D7",x"52",x"9D",x"AC",x"24",x"22",x"D6",x"42",x"D0",x"43",x"D7",x"42",x"80",x"30",x"34",
    x"02",x"8D",x"DB",x"26",x"BC",x"C6",x"0A",x"DD",x"5A",x"BD",x"D2",x"F2",x"8D",x"D0",x"26",x"C0",
    x"35",x"04",x"DD",x"5A",x"BD",x"D2",x"B0",x"20",x"DA",x"81",x"2E",x"27",x"31",x"81",x"21",x"27",
    x"39",x"81",x"45",x"26",x"39",x"9D",x"E9",x"8D",x"0E",x"D7",x"45",x"9D",x"AC",x"25",x"4A",x"0D",
    x"45",x"27",x"2B",x"00",x"44",x"20",x"27",x"9D",x"AC",x"5F",x"81",x"2D",x"27",x"0E",x"81",x"C8",
    x"27",x"0A",x"81",x"2B",x"27",x"07",x"81",x"C7",x"27",x"03",x"0E",x"CA",x"53",x"39",x"03",x"43",
    x"27",x"0C",x"8D",x"8A",x"26",x"9D",x"8D",x"6E",x"20",x"99",x"9D",x"E9",x"9D",x"AC",x"96",x"44",
    x"90",x"42",x"97",x"44",x"27",x"0E",x"2A",x"05",x"BD",x"DB",x"2A",x"20",x"07",x"BD",x"D4",x"B1",
    x"0A",x"44",x"26",x"F9",x"96",x"52",x"2B",x"17",x"39",x"C6",x"0A",x"D1",x"44",x"23",x"0A",x"34",
    x"02",x"96",x"44",x"3D",x"EB",x"E0",x"C0",x"30",x"8C",x"C6",x"32",x"D7",x"44",x"20",x"9C",x"9D",
    x"C5",x"2B",x"51",x"0D",x"4C",x"27",x"02",x"03",x"50",x"39",x"8D",x"1F",x"7E",x"D3",x"96",x"9D",
    x"C5",x"2A",x"F9",x"DC",x"4E",x"93",x"5A",x"29",x"F1",x"DD",x"4E",x"39",x"9D",x"C5",x"2A",x"08",
    x"DC",x"4E",x"D3",x"5A",x"28",x"F3",x"8D",x"03",x"7E",x"D3",x"9B",x"8D",x"09",x"DC",x"5A",x"34",
    x"06",x"BD",x"D6",x"80",x"20",x"04",x"DC",x"4E",x"34",x"06",x"8D",x"15",x"CC",x"04",x"90",x"DD",
    x"4B",x"EC",x"E1",x"27",x"0C",x"2A",x"05",x"03",x"50",x"BD",x"FF",x"3B",x"DD",x"4D",x"7E",x"D3",
    x"EF",x"7E",x"D4",x"54",x"8D",x"5D",x"29",x"43",x"39",x"8D",x"D0",x"7E",x"D4",x"B7",x"9D",x"C5",
    x"2A",x"F9",x"8D",x"3B",x"27",x"B3",x"DC",x"5A",x"27",x"AF",x"4D",x"26",x"1C",x"96",x"4E",x"3D",
    x"4D",x"26",x"E6",x"5D",x"2B",x"E3",x"6F",x"E2",x"34",x"04",x"96",x"4F",x"D6",x"5B",x"3D",x"E3",
    x"E1",x"29",x"D6",x"2B",x"0C",x"DD",x"4E",x"20",x"59",x"D6",x"4E",x"26",x"CC",x"D6",x"4F",x"20",
    x"DE",x"10",x"83",x"80",x"00",x"26",x"C2",x"0D",x"5D",x"2B",x"BD",x"4F",x"5F",x"20",x"97",x"96",
    x"4E",x"98",x"5A",x"97",x"5D",x"96",x"5A",x"2A",x"06",x"4F",x"5F",x"93",x"5A",x"DD",x"5A",x"DC",
    x"4E",x"2A",x"06",x"4F",x"5F",x"93",x"4E",x"DD",x"4E",x"39",x"DC",x"5A",x"10",x"27",x"01",x"91",
    x"8D",x"DD",x"86",x"10",x"97",x"4D",x"4F",x"5F",x"20",x"0C",x"93",x"5A",x"24",x"06",x"D3",x"5A",
    x"1C",x"FE",x"20",x"02",x"1A",x"01",x"DD",x"58",x"09",x"4F",x"09",x"4E",x"59",x"49",x"0A",x"4D",
    x"2A",x"E8",x"0D",x"5D",x"2B",x"CD",x"39",x"96",x"4E",x"34",x"02",x"8D",x"CD",x"DC",x"58",x"DD",
    x"4E",x"6D",x"E0",x"20",x"EF",x"EC",x"81",x"97",x"58",x"D7",x"5C",x"CA",x"80",x"D7",x"59",x"EC",
    x"81",x"DD",x"5A",x"39",x"8D",x"EF",x"03",x"50",x"8C",x"8D",x"EA",x"96",x"58",x"27",x"F4",x"D6",
    x"4C",x"10",x"27",x"02",x"CD",x"0F",x"51",x"D6",x"5C",x"D8",x"50",x"D7",x"5D",x"8E",x"21",x"58",
    x"D6",x"58",x"D0",x"4C",x"27",x"11",x"25",x"0A",x"97",x"4C",x"96",x"5C",x"97",x"50",x"8E",x"21",
    x"4C",x"50",x"BD",x"D4",x"5F",x"97",x"51",x"5F",x"DA",x"5D",x"2A",x"0D",x"63",x"01",x"63",x"02",
    x"63",x"03",x"96",x"51",x"43",x"89",x"00",x"97",x"51",x"DC",x"4E",x"D9",x"5B",x"99",x"5A",x"DD",
    x"4E",x"96",x"4D",x"99",x"59",x"97",x"4D",x"D6",x"5D",x"2A",x"41",x"25",x"02",x"8D",x"52",x"96",
    x"4D",x"2B",x"32",x"5F",x"D7",x"02",x"96",x"4D",x"26",x"14",x"DC",x"4E",x"DD",x"4D",x"96",x"51",
    x"97",x"4F",x"0A",x"02",x"0F",x"51",x"D6",x"02",x"C1",x"FC",x"26",x"EA",x"20",x"46",x"58",x"58",
    x"58",x"4D",x"20",x"09",x"5A",x"08",x"51",x"09",x"4F",x"09",x"4E",x"09",x"4D",x"2A",x"F5",x"DB",
    x"4C",x"D7",x"4C",x"24",x"2F",x"4F",x"08",x"51",x"97",x"51",x"20",x"0E",x"24",x"F7",x"0C",x"4C",
    x"10",x"27",x"00",x"AA",x"06",x"4D",x"06",x"4E",x"06",x"4F",x"24",x"04",x"8D",x"0B",x"27",x"EE",
    x"39",x"03",x"50",x"03",x"4D",x"03",x"4E",x"03",x"4F",x"0C",x"4F",x"26",x"06",x"0C",x"4E",x"26",
    x"02",x"0C",x"4D",x"39",x"0F",x"4E",x"0F",x"4F",x"4F",x"5F",x"DD",x"4C",x"DD",x"50",x"39",x"C1",
    x"F8",x"2F",x"1A",x"4F",x"07",x"56",x"66",x"01",x"20",x"1F",x"8E",x"21",x"0D",x"A6",x"03",x"34",
    x"04",x"97",x"51",x"EC",x"01",x"ED",x"02",x"96",x"56",x"A7",x"01",x"35",x"04",x"CB",x"08",x"2F",
    x"EC",x"96",x"51",x"C0",x"08",x"27",x"0A",x"67",x"01",x"66",x"02",x"66",x"03",x"46",x"5C",x"26",
    x"F6",x"39",x"4F",x"5F",x"DD",x"0E",x"DD",x"0F",x"D6",x"4F",x"8D",x"49",x"D6",x"51",x"D7",x"A5",
    x"D6",x"4E",x"8D",x"41",x"D6",x"51",x"D7",x"A4",x"D6",x"4D",x"8D",x"3B",x"D6",x"51",x"D7",x"A3",
    x"39",x"8E",x"DC",x"7D",x"BD",x"D3",x"85",x"8D",x"51",x"27",x"99",x"4D",x"27",x"96",x"34",x"04",
    x"8D",x"D0",x"BD",x"DB",x"A1",x"86",x"80",x"97",x"4C",x"BD",x"D3",x"EF",x"4F",x"D6",x"58",x"EB",
    x"E0",x"89",x"00",x"DB",x"4C",x"D7",x"4C",x"89",x"00",x"27",x"DE",x"4A",x"27",x"36",x"C6",x"06",
    x"8C",x"C6",x"0B",x"0E",x"FB",x"27",x"83",x"43",x"56",x"27",x"A6",x"34",x"04",x"24",x"0E",x"DC",
    x"0F",x"DB",x"5B",x"99",x"5A",x"DD",x"0F",x"96",x"0E",x"99",x"59",x"97",x"0E",x"06",x"0E",x"06",
    x"0F",x"06",x"10",x"06",x"51",x"5F",x"EA",x"E0",x"20",x"DE",x"96",x"5C",x"98",x"50",x"97",x"50",
    x"96",x"58",x"D6",x"4C",x"39",x"56",x"56",x"56",x"D7",x"51",x"20",x"A6",x"9D",x"C5",x"2A",x"08",
    x"BD",x"D2",x"BB",x"20",x"03",x"BD",x"D3",x"85",x"8D",x"E0",x"27",x"B5",x"4D",x"27",x"AA",x"50",
    x"5C",x"34",x"04",x"8E",x"21",x"0E",x"CC",x"03",x"01",x"97",x"02",x"8D",x"38",x"26",x"01",x"43",
    x"1F",x"A8",x"59",x"24",x"0E",x"0D",x"02",x"27",x"CC",x"E7",x"80",x"C6",x"01",x"0A",x"02",x"26",
    x"02",x"C6",x"40",x"34",x"04",x"1F",x"8A",x"24",x"0E",x"DC",x"5A",x"D0",x"4F",x"92",x"4E",x"DD",
    x"5A",x"96",x"59",x"92",x"4D",x"97",x"59",x"08",x"5B",x"09",x"5A",x"09",x"59",x"35",x"04",x"25",
    x"CF",x"2B",x"C8",x"20",x"CB",x"34",x"04",x"DC",x"4D",x"93",x"59",x"26",x"04",x"96",x"4F",x"90",
    x"5B",x"35",x"84",x"9D",x"D1",x"2A",x"0B",x"DC",x"4E",x"26",x"0D",x"4F",x"5F",x"39",x"CC",x"00",
    x"01",x"39",x"D6",x"4C",x"27",x"F5",x"D6",x"50",x"2A",x"F4",x"CC",x"FF",x"FF",x"39",x"8D",x"E3",
    x"2A",x"EB",x"7E",x"D2",x"8F",x"D6",x"5A",x"96",x"4E",x"98",x"5A",x"2B",x"07",x"DC",x"5A",x"93",
    x"4E",x"27",x"D8",x"56",x"5D",x"20",x"E1",x"9D",x"C5",x"2B",x"EA",x"D6",x"5C",x"96",x"50",x"98",
    x"5C",x"2B",x"F1",x"96",x"4C",x"91",x"58",x"26",x"05",x"4D",x"27",x"BF",x"8D",x"A7",x"8D",x"E1",
    x"27",x"35",x"0D",x"5C",x"2B",x"31",x"7E",x"FF",x"3B",x"8D",x"A8",x"1D",x"DD",x"4E",x"20",x"71",
    x"9D",x"C5",x"2B",x"23",x"8D",x"9D",x"2A",x"20",x"03",x"50",x"8D",x"1C",x"20",x"B4",x"D6",x"4C",
    x"10",x"27",x"FE",x"60",x"C0",x"98",x"96",x"50",x"2A",x"05",x"03",x"56",x"BD",x"D4",x"43",x"8E",
    x"21",x"4C",x"BD",x"D4",x"5F",x"0F",x"56",x"39",x"D6",x"4C",x"8D",x"4C",x"2B",x"F9",x"C1",x"98",
    x"24",x"F5",x"8D",x"DA",x"D7",x"51",x"96",x"50",x"D7",x"50",x"80",x"80",x"86",x"98",x"97",x"4C",
    x"96",x"4F",x"97",x"00",x"7E",x"D3",x"EB",x"8D",x"2F",x"2B",x"2A",x"D6",x"4C",x"27",x"AC",x"C1",
    x"90",x"25",x"03",x"7E",x"D4",x"DE",x"96",x"50",x"34",x"02",x"0F",x"50",x"8D",x"B0",x"4D",x"2A",
    x"09",x"DC",x"4E",x"C3",x"00",x"01",x"29",x"EB",x"DD",x"4E",x"A6",x"E0",x"2A",x"03",x"BD",x"D3",
    x"43",x"86",x"02",x"97",x"4B",x"DC",x"4E",x"39",x"9D",x"C5",x"26",x"FB",x"C6",x"0D",x"0E",x"FB",
    x"9D",x"C5",x"26",x"F8",x"39",x"9D",x"C7",x"27",x"F7",x"2B",x"BC",x"8D",x"EB",x"29",x"E8",x"7E",
    x"D2",x"C6",x"96",x"5C",x"5F",x"DD",x"50",x"DC",x"58",x"DD",x"4C",x"DC",x"5A",x"DD",x"4E",x"39",
    x"96",x"50",x"97",x"5C",x"DC",x"4E",x"DD",x"5A",x"DC",x"4C",x"DD",x"58",x"39",x"9D",x"C5",x"2B",
    x"15",x"EC",x"02",x"DD",x"4E",x"0F",x"51",x"EC",x"84",x"97",x"4C",x"10",x"27",x"FD",x"B5",x"D7",
    x"50",x"CA",x"80",x"D7",x"4D",x"39",x"EC",x"84",x"DD",x"4E",x"39",x"9D",x"E9",x"8D",x"D1",x"8E",
    x"DC",x"79",x"8D",x"D9",x"96",x"4C",x"27",x"7C",x"96",x"58",x"26",x"07",x"0D",x"50",x"2A",x"71",
    x"7E",x"D4",x"E1",x"8E",x"21",x"46",x"BD",x"D7",x"F3",x"5F",x"96",x"5C",x"2A",x"0F",x"BD",x"D6",
    x"08",x"8E",x"21",x"46",x"BD",x"DC",x"00",x"26",x"04",x"03",x"5C",x"D6",x"00",x"34",x"04",x"8D",
    x"91",x"8D",x"0E",x"8E",x"21",x"46",x"8D",x"47",x"8D",x"4A",x"66",x"E0",x"10",x"25",x"FB",x"9F",
    x"39",x"9D",x"E9",x"BD",x"D5",x"83",x"10",x"2F",x"4A",x"FC",x"8E",x"DC",x"44",x"96",x"4C",x"80",
    x"80",x"34",x"02",x"86",x"80",x"97",x"4C",x"8D",x"69",x"8E",x"DC",x"48",x"BD",x"D5",x"25",x"8E",
    x"DC",x"33",x"BD",x"D3",x"94",x"8E",x"DC",x"37",x"8D",x"62",x"8E",x"DC",x"4C",x"8D",x"53",x"8D",
    x"70",x"35",x"04",x"1D",x"BD",x"D2",x"C8",x"8E",x"21",x"3E",x"8D",x"46",x"8E",x"DC",x"50",x"20",
    x"56",x"7E",x"D4",x"54",x"8D",x"59",x"8E",x"DC",x"54",x"8D",x"4C",x"96",x"4C",x"81",x"88",x"24",
    x"34",x"BD",x"D6",x"08",x"96",x"00",x"8B",x"81",x"27",x"2B",x"34",x"02",x"8E",x"DC",x"33",x"8D",
    x"D9",x"8E",x"21",x"3E",x"BD",x"D3",x"94",x"BD",x"D2",x"93",x"10",x"8E",x"DC",x"58",x"8D",x"36",
    x"96",x"4C",x"80",x"80",x"AB",x"E0",x"29",x"11",x"27",x"C7",x"97",x"4C",x"0F",x"50",x"39",x"8E",
    x"DC",x"79",x"7E",x"D3",x"99",x"96",x"50",x"2B",x"B8",x"7E",x"D4",x"DE",x"1F",x"12",x"8D",x"11",
    x"8D",x"05",x"8D",x"12",x"8E",x"21",x"3E",x"7E",x"D4",x"B4",x"8E",x"21",x"42",x"20",x"68",x"9D",
    x"E9",x"8E",x"21",x"3E",x"20",x"61",x"8D",x"F2",x"E6",x"A0",x"D7",x"52",x"1F",x"21",x"8D",x"E7",
    x"31",x"24",x"1F",x"21",x"8D",x"CC",x"8E",x"21",x"42",x"0A",x"52",x"26",x"F1",x"39",x"9D",x"E9",
    x"8E",x"DC",x"12",x"8D",x"BD",x"9D",x"E9",x"96",x"4C",x"81",x"77",x"25",x"F0",x"8E",x"DC",x"16",
    x"8D",x"C5",x"BD",x"D6",x"80",x"BD",x"D6",x"08",x"BD",x"D3",x"96",x"8E",x"DC",x"1A",x"BD",x"D3",
    x"94",x"96",x"50",x"34",x"02",x"2A",x"06",x"8D",x"96",x"96",x"50",x"2B",x"03",x"BD",x"D2",x"93",
    x"8E",x"DC",x"1A",x"8D",x"8D",x"A6",x"E0",x"2A",x"03",x"BD",x"D2",x"93",x"8E",x"DC",x"1E",x"20",
    x"8B",x"9E",x"3B",x"9D",x"C5",x"28",x"0F",x"96",x"4C",x"D6",x"50",x"CA",x"7F",x"D4",x"4D",x"ED",
    x"84",x"DC",x"4E",x"ED",x"02",x"39",x"DC",x"4E",x"ED",x"84",x"39",x"BD",x"C7",x"E3",x"8D",x"A5",
    x"8E",x"21",x"46",x"BD",x"D7",x"F3",x"BD",x"C7",x"FB",x"8D",x"93",x"8E",x"21",x"46",x"7E",x"D5",
    x"25",x"4A",x"4A",x"4A",x"2F",x"02",x"1A",x"02",x"39",x"0D",x"B4",x"26",x"02",x"0A",x"B3",x"0A",
    x"B4",x"39",x"20",x"69",x"6E",x"20",x"00",x"8E",x"D8",x"31",x"8D",x"06",x"DC",x"24",x"8D",x"05",
    x"8D",x"10",x"7E",x"CE",x"2C",x"DD",x"4E",x"BD",x"D4",x"58",x"CC",x"04",x"98",x"DD",x"4B",x"7E",
    x"D3",x"EF",x"0F",x"78",x"8E",x"25",x"56",x"9F",x"5E",x"C6",x"20",x"96",x"78",x"85",x"08",x"27",
    x"02",x"C6",x"2B",x"34",x"04",x"BD",x"D5",x"83",x"35",x"02",x"34",x"04",x"2A",x"05",x"BD",x"D2",
    x"8F",x"86",x"2D",x"BD",x"D9",x"F8",x"9E",x"5E",x"C6",x"30",x"E7",x"80",x"96",x"78",x"35",x"04",
    x"10",x"2B",x"01",x"7E",x"5D",x"26",x"05",x"6F",x"84",x"30",x"1E",x"39",x"0F",x"42",x"9D",x"C5",
    x"2A",x"64",x"BD",x"D9",x"C1",x"8E",x"25",x"56",x"E6",x"84",x"86",x"20",x"34",x"04",x"D6",x"78",
    x"C5",x"20",x"35",x"04",x"27",x"08",x"86",x"2A",x"C1",x"20",x"26",x"02",x"1F",x"89",x"34",x"04",
    x"A7",x"80",x"E6",x"84",x"27",x"10",x"C1",x"45",x"27",x"0C",x"C1",x"30",x"27",x"F2",x"C1",x"2C",
    x"27",x"EE",x"C1",x"2E",x"26",x"04",x"86",x"30",x"A7",x"82",x"35",x"04",x"E7",x"82",x"39",x"4A",
    x"97",x"44",x"BD",x"C7",x"E3",x"8D",x"37",x"BD",x"C7",x"FB",x"D6",x"44",x"53",x"96",x"42",x"34",
    x"04",x"A1",x"E0",x"25",x"5F",x"34",x"04",x"8E",x"25",x"57",x"9F",x"5E",x"BD",x"D9",x"EA",x"A6",
    x"E0",x"BD",x"DA",x"73",x"20",x"11",x"8D",x"50",x"96",x"44",x"C6",x"02",x"D7",x"42",x"8B",x"06",
    x"2B",x"CD",x"81",x"06",x"2E",x"05",x"4C",x"97",x"42",x"86",x"01",x"4A",x"97",x"44",x"8D",x"6B",
    x"C6",x"FF",x"5C",x"A6",x"82",x"81",x"30",x"27",x"F9",x"81",x"2E",x"27",x"02",x"30",x"01",x"D7",
    x"42",x"6F",x"84",x"D6",x"44",x"27",x"1D",x"86",x"2B",x"5D",x"2A",x"03",x"86",x"2D",x"50",x"A7",
    x"01",x"86",x"45",x"A7",x"81",x"86",x"2F",x"4C",x"C0",x"0A",x"24",x"FB",x"CB",x"3A",x"ED",x"81",
    x"6F",x"84",x"9F",x"5E",x"8E",x"25",x"56",x"39",x"4F",x"97",x"44",x"D6",x"4C",x"8E",x"DB",x"84",
    x"E1",x"80",x"22",x"09",x"BD",x"D4",x"B4",x"86",x"FA",x"9B",x"44",x"20",x"EC",x"8E",x"DB",x"8D",
    x"BD",x"DC",x"00",x"23",x"07",x"BD",x"DB",x"95",x"0C",x"44",x"20",x"F1",x"8E",x"DB",x"89",x"BD",
    x"DC",x"00",x"22",x"D3",x"BD",x"D4",x"B1",x"0A",x"44",x"20",x"F1",x"BD",x"D7",x"6F",x"BD",x"D5",
    x"EE",x"8E",x"DB",x"74",x"C6",x"80",x"8D",x"5E",x"4F",x"8D",x"0D",x"28",x"FB",x"8D",x"1F",x"8C",
    x"DB",x"7A",x"26",x"F2",x"30",x"02",x"20",x"2C",x"96",x"4F",x"A9",x"02",x"97",x"4F",x"96",x"4E",
    x"A9",x"01",x"97",x"4E",x"96",x"4D",x"A9",x"84",x"97",x"4D",x"5C",x"56",x"59",x"39",x"30",x"03",
    x"24",x"03",x"C0",x"0B",x"50",x"CB",x"2F",x"1F",x"98",x"84",x"7F",x"8D",x"3B",x"53",x"C4",x"80",
    x"39",x"8E",x"DB",x"7A",x"8D",x"20",x"86",x"2F",x"34",x"02",x"DC",x"4E",x"6C",x"E4",x"DD",x"4E",
    x"A3",x"84",x"24",x"F8",x"30",x"02",x"A6",x"E0",x"8D",x"1E",x"8C",x"DB",x"84",x"26",x"E5",x"8D",
    x"05",x"9E",x"5E",x"6F",x"84",x"39",x"0A",x"42",x"26",x"FB",x"86",x"2E",x"34",x"10",x"8D",x"08",
    x"9E",x"5E",x"30",x"1F",x"9F",x"37",x"35",x"90",x"34",x"10",x"9E",x"5E",x"A7",x"80",x"9F",x"5E",
    x"35",x"90",x"9F",x"5E",x"9D",x"C5",x"10",x"2A",x"00",x"90",x"96",x"78",x"46",x"10",x"25",x"01",
    x"1C",x"86",x"06",x"97",x"42",x"96",x"77",x"80",x"05",x"8D",x"58",x"8D",x"A4",x"96",x"76",x"26",
    x"04",x"30",x"1F",x"9F",x"5E",x"4A",x"8D",x"4B",x"BD",x"D8",x"95",x"4F",x"8D",x"CA",x"8E",x"25",
    x"55",x"30",x"01",x"9F",x"0A",x"96",x"38",x"90",x"0B",x"90",x"77",x"27",x"A8",x"A6",x"84",x"81",
    x"20",x"27",x"EE",x"81",x"2A",x"27",x"EA",x"4F",x"34",x"02",x"A6",x"80",x"81",x"2D",x"27",x"F8",
    x"81",x"2B",x"27",x"F4",x"81",x"30",x"26",x"0E",x"A6",x"01",x"9D",x"B9",x"24",x"08",x"35",x"02",
    x"A7",x"82",x"26",x"FA",x"20",x"CB",x"A6",x"E0",x"26",x"FC",x"9E",x"0A",x"86",x"25",x"A7",x"82",
    x"39",x"8D",x"1E",x"4A",x"2A",x"FB",x"39",x"96",x"44",x"34",x"04",x"AB",x"E0",x"4C",x"97",x"42",
    x"39",x"34",x"02",x"BD",x"D9",x"E6",x"35",x"02",x"4A",x"2B",x"05",x"8D",x"04",x"4D",x"26",x"F1",
    x"39",x"34",x"02",x"86",x"30",x"BD",x"D9",x"F8",x"35",x"82",x"96",x"78",x"46",x"10",x"25",x"00",
    x"8F",x"8E",x"DB",x"91",x"BD",x"DC",x"00",x"25",x"05",x"BD",x"D8",x"52",x"20",x"BE",x"C6",x"06",
    x"96",x"4C",x"97",x"44",x"27",x"05",x"BD",x"D9",x"48",x"C6",x"06",x"96",x"44",x"2B",x"25",x"40",
    x"9B",x"77",x"34",x"04",x"A0",x"E0",x"8D",x"AB",x"8D",x"AD",x"BD",x"D9",x"7B",x"96",x"44",x"8D",
    x"B7",x"96",x"44",x"BD",x"D9",x"E6",x"9E",x"5E",x"7E",x"DA",x"1D",x"34",x"04",x"A0",x"E0",x"90",
    x"44",x"7E",x"DA",x"73",x"96",x"76",x"27",x"01",x"4A",x"9B",x"44",x"2B",x"01",x"4F",x"34",x"06",
    x"8D",x"38",x"96",x"44",x"A0",x"E0",x"97",x"44",x"AB",x"E4",x"35",x"04",x"2B",x"09",x"96",x"77",
    x"8D",x"D9",x"BD",x"DA",x"77",x"20",x"0C",x"96",x"77",x"8D",x"D6",x"BD",x"D9",x"EA",x"4F",x"8D",
    x"CA",x"0F",x"42",x"BD",x"D9",x"7B",x"96",x"76",x"26",x"04",x"9E",x"37",x"9F",x"5E",x"9B",x"44",
    x"7E",x"DA",x"25",x"34",x"02",x"8D",x"6E",x"35",x"02",x"4C",x"2B",x"F7",x"39",x"BD",x"D2",x"C6",
    x"96",x"4C",x"34",x"02",x"27",x"03",x"BD",x"D9",x"48",x"96",x"76",x"27",x"01",x"4A",x"9B",x"77",
    x"4A",x"80",x"06",x"34",x"02",x"8D",x"E3",x"A6",x"E4",x"2B",x"01",x"4F",x"40",x"9B",x"77",x"97",
    x"42",x"BD",x"D9",x"7B",x"35",x"02",x"BD",x"DA",x"88",x"9E",x"5E",x"96",x"76",x"26",x"02",x"30",
    x"1F",x"E6",x"E0",x"27",x"07",x"D6",x"44",x"CB",x"06",x"D0",x"77",x"5C",x"BD",x"D9",x"27",x"9E",
    x"5E",x"7E",x"DA",x"28",x"FE",x"79",x"60",x"00",x"27",x"10",x"27",x"10",x"03",x"E8",x"00",x"64",
    x"00",x"0A",x"00",x"01",x"80",x"94",x"74",x"24",x"00",x"91",x"43",x"4F",x"F8",x"94",x"74",x"23",
    x"F7",x"B6",x"0E",x"1B",x"C9",x"BD",x"D6",x"80",x"8E",x"DC",x"7D",x"BD",x"D6",x"8D",x"7E",x"D5",
    x"28",x"DC",x"0E",x"DD",x"4D",x"96",x"10",x"97",x"4F",x"39",x"86",x"04",x"97",x"4B",x"8E",x"DC",
    x"33",x"BD",x"D6",x"8D",x"20",x"0B",x"9D",x"B2",x"81",x"28",x"26",x"EE",x"BD",x"C7",x"29",x"9D",
    x"E9",x"10",x"8E",x"24",x"27",x"BD",x"D5",x"83",x"2B",x"0A",x"27",x"23",x"EC",x"21",x"DD",x"4D",
    x"A6",x"23",x"97",x"4F",x"CC",x"40",x"E6",x"DD",x"59",x"86",x"4D",x"97",x"5B",x"BD",x"D4",x"92",
    x"DC",x"A4",x"C3",x"B0",x"65",x"ED",x"22",x"D6",x"A3",x"C9",x"05",x"96",x"0F",x"ED",x"A4",x"EC",
    x"A4",x"97",x"51",x"86",x"80",x"DD",x"4C",x"EC",x"22",x"DD",x"4E",x"0F",x"50",x"7E",x"D3",x"EF",
    x"34",x"02",x"DC",x"4C",x"C4",x"7F",x"10",x"A3",x"84",x"26",x"05",x"DC",x"4E",x"10",x"A3",x"02",
    x"35",x"82",x"81",x"49",x"0F",x"DB",x"7E",x"22",x"F9",x"83",x"7F",x"00",x"00",x"00",x"04",x"86",
    x"1E",x"D7",x"BA",x"87",x"99",x"26",x"64",x"87",x"23",x"34",x"58",x"86",x"A5",x"5D",x"E0",x"83",
    x"49",x"0F",x"DA",x"81",x"00",x"00",x"00",x"02",x"80",x"19",x"56",x"AA",x"80",x"76",x"22",x"F1",
    x"82",x"38",x"AA",x"45",x"80",x"35",x"04",x"F3",x"81",x"35",x"04",x"F3",x"80",x"80",x"00",x"00",
    x"80",x"31",x"72",x"18",x"81",x"38",x"AA",x"3B",x"07",x"74",x"94",x"2E",x"40",x"77",x"2E",x"4F",
    x"70",x"7A",x"88",x"02",x"6E",x"7C",x"2A",x"A0",x"E6",x"7E",x"AA",x"AA",x"50",x"7F",x"7F",x"FF",
    x"FF",x"81",x"80",x"00",x"00",x"81",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"84",x"20",x"00",
    x"00",x"9D",x"AC",x"C6",x"A1",x"9D",x"E0",x"8D",x"1E",x"8D",x"70",x"0F",x"79",x"9D",x"F0",x"9F",
    x"3B",x"9D",x"D6",x"8E",x"24",x"51",x"4F",x"BD",x"CB",x"71",x"7E",x"C6",x"7C",x"9D",x"AC",x"D6",
    x"4A",x"10",x"26",x"F1",x"97",x"39",x"C6",x"5F",x"D7",x"4A",x"C6",x"0C",x"9E",x"24",x"30",x"01",
    x"27",x"56",x"81",x"3B",x"26",x"02",x"9D",x"AC",x"81",x"23",x"26",x"0A",x"BD",x"E1",x"D0",x"9D",
    x"C2",x"BD",x"E4",x"19",x"9D",x"B2",x"81",x"22",x"26",x"D5",x"BD",x"C6",x"E1",x"BD",x"CE",x"2F",
    x"9D",x"B2",x"81",x"3B",x"27",x"C7",x"0E",x"C2",x"9E",x"2E",x"9F",x"24",x"0E",x"F9",x"9F",x"B3",
    x"BD",x"C5",x"7D",x"6D",x"80",x"26",x"0A",x"C6",x"04",x"EE",x"81",x"27",x"1B",x"EC",x"81",x"DD",
    x"2E",x"9F",x"B3",x"9D",x"B2",x"81",x"83",x"26",x"E7",x"20",x"6E",x"BD",x"EC",x"CF",x"10",x"25",
    x"E7",x"AD",x"C6",x"36",x"0D",x"7A",x"27",x"9D",x"0E",x"FB",x"9D",x"AC",x"81",x"B8",x"10",x"27",
    x"0B",x"A8",x"8D",x"92",x"4F",x"BD",x"E3",x"B6",x"2B",x"04",x"8D",x"DF",x"86",x"2C",x"8E",x"24",
    x"51",x"A7",x"84",x"20",x"19",x"C6",x"3A",x"BD",x"E3",x"B6",x"26",x"DC",x"96",x"04",x"26",x"A8",
    x"8E",x"DD",x"D1",x"BD",x"CE",x"2C",x"9E",x"2C",x"9F",x"B3",x"39",x"9E",x"30",x"86",x"4F",x"97",
    x"04",x"9F",x"32",x"8C",x"9D",x"C2",x"9D",x"F0",x"9F",x"3B",x"9E",x"B3",x"9F",x"28",x"9E",x"32",
    x"A6",x"84",x"9D",x"B9",x"26",x"11",x"96",x"04",x"26",x"84",x"BD",x"E3",x"B6",x"27",x"C6",x"2A",
    x"04",x"BD",x"22",x"6C",x"8C",x"8D",x"94",x"9F",x"B3",x"9D",x"C5",x"27",x"43",x"9E",x"B3",x"9D",
    x"AC",x"DE",x"B3",x"34",x"40",x"9F",x"B3",x"96",x"4B",x"34",x"02",x"BD",x"D1",x"E3",x"35",x"02",
    x"BD",x"D6",x"65",x"9E",x"B3",x"AC",x"E1",x"27",x"D4",x"BD",x"D7",x"F1",x"9D",x"B2",x"27",x"04",
    x"81",x"2C",x"26",x"91",x"9E",x"B3",x"9F",x"32",x"9E",x"28",x"9F",x"B3",x"9D",x"B2",x"26",x"A4",
    x"9E",x"32",x"D6",x"04",x"27",x"03",x"9F",x"30",x"39",x"A6",x"84",x"26",x"83",x"0F",x"79",x"39",
    x"4F",x"5F",x"9D",x"F3",x"0D",x"8F",x"26",x"0F",x"9D",x"AC",x"9E",x"B3",x"1F",x"89",x"81",x"22",
    x"27",x"05",x"30",x"1F",x"CC",x"3A",x"2C",x"BD",x"CB",x"73",x"BD",x"C6",x"E6",x"BD",x"C6",x"7C",
    x"20",x"BA",x"3F",x"52",x"65",x"64",x"6F",x"0D",x"0A",x"00",x"BD",x"E1",x"07",x"30",x"04",x"10",
    x"8E",x"24",x"52",x"EC",x"80",x"4D",x"27",x"4C",x"2B",x"0F",x"81",x"3A",x"26",x"08",x"C1",x"8F",
    x"27",x"F1",x"C1",x"8D",x"27",x"ED",x"8D",x"32",x"8C",x"8D",x"02",x"20",x"E6",x"CE",x"21",x"F7",
    x"81",x"FF",x"26",x"06",x"1F",x"98",x"33",x"45",x"30",x"01",x"84",x"7F",x"33",x"4A",x"A0",x"C4",
    x"2A",x"FA",x"AB",x"C4",x"EE",x"41",x"4A",x"2B",x"06",x"6D",x"C0",x"2A",x"FC",x"20",x"F7",x"A6",
    x"C4",x"84",x"7F",x"8D",x"05",x"6D",x"C0",x"2A",x"F6",x"39",x"10",x"8C",x"25",x"51",x"24",x"04",
    x"A7",x"A0",x"6F",x"A4",x"39",x"86",x"AB",x"A7",x"C0",x"39",x"CE",x"24",x"51",x"A6",x"80",x"A7",
    x"C0",x"27",x"18",x"9D",x"B9",x"25",x"F6",x"33",x"5F",x"10",x"8E",x"DF",x"0C",x"A1",x"A1",x"25",
    x"FC",x"26",x"2D",x"E6",x"A2",x"1F",x"52",x"AD",x"A5",x"26",x"E2",x"5F",x"ED",x"C1",x"1F",x"30",
    x"83",x"24",x"4F",x"8E",x"24",x"50",x"9F",x"B3",x"39",x"CC",x"3A",x"8D",x"ED",x"C1",x"4F",x"8C",
    x"A7",x"C0",x"97",x"3F",x"A6",x"80",x"A7",x"C0",x"27",x"05",x"91",x"3F",x"26",x"F6",x"43",x"39",
    x"30",x"1F",x"34",x"50",x"0F",x"3E",x"CE",x"21",x"F7",x"0F",x"3F",x"33",x"4A",x"E6",x"C4",x"27",
    x"36",x"10",x"AE",x"41",x"AE",x"E4",x"A6",x"80",x"8D",x"5F",x"A0",x"A0",x"27",x"F8",x"81",x"80",
    x"26",x"45",x"35",x"60",x"9A",x"3F",x"D6",x"3E",x"26",x"06",x"81",x"8F",x"26",x"04",x"C6",x"3A",
    x"E7",x"C0",x"A7",x"C0",x"5C",x"27",x"86",x"8D",x"02",x"20",x"9E",x"81",x"8C",x"27",x"AF",x"81",
    x"83",x"26",x"BB",x"86",x"00",x"20",x"AB",x"CE",x"21",x"FC",x"03",x"3E",x"26",x"BB",x"35",x"50",
    x"A6",x"80",x"8D",x"20",x"24",x"DC",x"A7",x"C0",x"27",x"81",x"A6",x"80",x"8D",x"16",x"25",x"F6",
    x"9D",x"B9",x"25",x"F2",x"7E",x"DE",x"3F",x"0C",x"3F",x"5A",x"27",x"9F",x"31",x"3F",x"A6",x"A0",
    x"2A",x"FC",x"20",x"A0",x"8D",x"03",x"7E",x"C8",x"A1",x"81",x"16",x"26",x"04",x"A6",x"01",x"30",
    x"02",x"81",x"61",x"25",x"06",x"81",x"7A",x"22",x"02",x"88",x"20",x"39",x"3F",x"DE",x"3A",x"E0",
    x"27",x"12",x"22",x"19",x"20",x"E0",x"00",x"96",x"24",x"4C",x"10",x"27",x"E5",x"94",x"0D",x"23",
    x"27",x"F8",x"C6",x"13",x"0E",x"FB",x"10",x"DF",x"72",x"BD",x"E4",x"79",x"9E",x"B3",x"9F",x"2C",
    x"A6",x"80",x"27",x"08",x"81",x"3A",x"27",x"22",x"0E",x"F9",x"03",x"23",x"4F",x"EC",x"81",x"27",
    x"D6",x"EC",x"80",x"DD",x"24",x"9F",x"B3",x"96",x"6E",x"27",x"0F",x"86",x"5B",x"BD",x"CE",x"46",
    x"96",x"24",x"BD",x"D8",x"3E",x"86",x"5D",x"BD",x"CE",x"46",x"9D",x"AC",x"8D",x"02",x"20",x"C6",
    x"27",x"A9",x"81",x"80",x"10",x"25",x"E7",x"07",x"81",x"B9",x"22",x"0B",x"BE",x"22",x"04",x"48",
    x"1F",x"89",x"3A",x"9D",x"AC",x"6E",x"94",x"81",x"FF",x"27",x"08",x"81",x"D5",x"23",x"B9",x"6E",
    x"9F",x"22",x"0E",x"9D",x"AC",x"81",x"A1",x"10",x"27",x"FD",x"7F",x"81",x"A4",x"10",x"27",x"07",
    x"19",x"7E",x"22",x"7B",x"96",x"8D",x"97",x"8E",x"8E",x"23",x"FA",x"6F",x"80",x"CC",x"20",x"08",
    x"A7",x"80",x"5A",x"26",x"FB",x"37",x"24",x"E7",x"84",x"10",x"AF",x"01",x"9D",x"B2",x"27",x"7C",
    x"BD",x"CB",x"F5",x"C1",x"02",x"25",x"31",x"86",x"3A",x"A1",x"01",x"27",x"34",x"C1",x"05",x"25",
    x"27",x"A1",x"04",x"26",x"23",x"34",x"14",x"C6",x"0F",x"D7",x"8E",x"CE",x"23",x"C8",x"D6",x"8E",
    x"58",x"EE",x"C5",x"27",x"15",x"AE",x"61",x"C6",x"04",x"A6",x"C0",x"A1",x"80",x"26",x"0B",x"5A",
    x"26",x"F7",x"35",x"14",x"30",x"05",x"C0",x"05",x"20",x"17",x"0A",x"8E",x"2A",x"DD",x"7E",x"E2",
    x"39",x"A6",x"81",x"80",x"30",x"25",x"29",x"81",x"09",x"22",x"25",x"8A",x"80",x"97",x"8E",x"C0",
    x"02",x"CE",x"24",x"06",x"5D",x"27",x"1E",x"A6",x"84",x"81",x"28",x"26",x"18",x"30",x"01",x"5A",
    x"27",x"0E",x"A6",x"80",x"81",x"29",x"27",x"0C",x"A7",x"C0",x"11",x"83",x"24",x"27",x"25",x"EF",
    x"C6",x"37",x"0E",x"FB",x"5A",x"6F",x"C4",x"CE",x"23",x"FB",x"5C",x"5A",x"27",x"3B",x"A6",x"80",
    x"81",x"2E",x"27",x"0D",x"11",x"83",x"24",x"03",x"27",x"E6",x"8D",x"21",x"7C",x"23",x"FA",x"20",
    x"EA",x"CE",x"24",x"06",x"86",x"20",x"A7",x"C2",x"11",x"83",x"24",x"03",x"26",x"F8",x"5A",x"27",
    x"18",x"A6",x"80",x"11",x"83",x"24",x"06",x"27",x"C7",x"8D",x"02",x"20",x"F1",x"A7",x"C0",x"10",
    x"8E",x"E4",x"59",x"A1",x"A0",x"27",x"B9",x"22",x"FA",x"39",x"81",x"22",x"26",x"1E",x"8D",x"06",
    x"27",x"1A",x"9D",x"C2",x"20",x"16",x"CE",x"E4",x"60",x"BD",x"DF",x"94",x"C6",x"11",x"D7",x"79",
    x"0F",x"91",x"0F",x"92",x"0F",x"96",x"0E",x"B2",x"9D",x"AC",x"26",x"5C",x"BD",x"CE",x"82",x"34",
    x"10",x"8D",x"74",x"03",x"92",x"03",x"96",x"0D",x"79",x"27",x"03",x"BD",x"E2",x"1F",x"35",x"50",
    x"7E",x"CE",x"4A",x"81",x"4D",x"10",x"27",x"00",x"AC",x"8D",x"CB",x"27",x"7C",x"9D",x"C2",x"81",
    x"41",x"27",x"D5",x"C6",x"50",x"9D",x"E0",x"26",x"2F",x"BD",x"E2",x"1F",x"8D",x"14",x"9C",x"15",
    x"27",x"4D",x"A6",x"84",x"90",x"4C",x"8D",x"12",x"8D",x"17",x"9B",x"4D",x"A7",x"80",x"8D",x"19",
    x"20",x"EC",x"CC",x"0B",x"0D",x"DD",x"4C",x"9E",x"13",x"39",x"CE",x"DC",x"37",x"D6",x"4C",x"20",
    x"05",x"CE",x"DC",x"1E",x"D6",x"4D",x"A8",x"C5",x"39",x"CC",x"0B",x"0D",x"0A",x"4C",x"26",x"02",
    x"97",x"4C",x"0A",x"4D",x"26",x"F2",x"D7",x"4D",x"39",x"9D",x"AC",x"CE",x"E4",x"66",x"BD",x"E0",
    x"79",x"9E",x"24",x"30",x"01",x"26",x"E1",x"0D",x"7F",x"27",x"DD",x"C6",x"3D",x"0E",x"FB",x"86",
    x"FE",x"8D",x"1D",x"8D",x"BD",x"9C",x"15",x"27",x"CF",x"A6",x"84",x"90",x"4D",x"8D",x"C2",x"8D",
    x"B9",x"9B",x"4C",x"A7",x"80",x"8D",x"C2",x"20",x"EC",x"8D",x"DC",x"BD",x"E2",x"1F",x"86",x"FF",
    x"9D",x"E3",x"DC",x"15",x"93",x"13",x"8D",x"17",x"9E",x"13",x"A6",x"80",x"9D",x"E3",x"9C",x"15",
    x"26",x"F8",x"20",x"52",x"9D",x"C2",x"BD",x"CC",x"BA",x"EE",x"E4",x"AF",x"E4",x"1F",x"35",x"9D",
    x"E3",x"1E",x"89",x"0E",x"E3",x"8D",x"A2",x"8D",x"EB",x"8D",x"E9",x"AC",x"62",x"10",x"25",x"40",
    x"95",x"8D",x"E1",x"9D",x"B2",x"26",x"50",x"86",x"02",x"97",x"91",x"BD",x"E2",x"1F",x"4F",x"8D",
    x"E2",x"EC",x"62",x"A3",x"64",x"C3",x"00",x"01",x"1F",x"02",x"8D",x"D3",x"EC",x"64",x"8D",x"CF",
    x"AE",x"64",x"A6",x"80",x"9D",x"E3",x"31",x"3F",x"26",x"F8",x"86",x"FF",x"8D",x"C5",x"4F",x"5F",
    x"8D",x"BD",x"35",x"36",x"8D",x"B9",x"D6",x"79",x"0F",x"79",x"8E",x"23",x"E8",x"A6",x"85",x"27",
    x"2C",x"10",x"2B",x"40",x"B8",x"34",x"14",x"84",x"30",x"97",x"90",x"E6",x"85",x"BD",x"E3",x"A2",
    x"AD",x"98",x"06",x"35",x"14",x"6F",x"85",x"39",x"27",x"0C",x"8D",x"14",x"8D",x"D8",x"9D",x"B2",
    x"27",x"0B",x"8D",x"0A",x"20",x"F6",x"C6",x"11",x"8D",x"CE",x"5A",x"2A",x"FB",x"39",x"9D",x"C2",
    x"9D",x"B2",x"81",x"23",x"26",x"02",x"9D",x"AC",x"9D",x"CD",x"BD",x"CC",x"B2",x"C1",x"10",x"22",
    x"04",x"D7",x"79",x"26",x"E8",x"C6",x"32",x"0E",x"FB",x"BD",x"CC",x"15",x"34",x"04",x"8D",x"DE",
    x"8E",x"23",x"E8",x"6D",x"85",x"26",x"3F",x"9D",x"C2",x"CE",x"E4",x"63",x"BD",x"DF",x"94",x"BD",
    x"22",x"6F",x"9D",x"B2",x"26",x"4C",x"CC",x"01",x"FF",x"DD",x"91",x"D7",x"96",x"35",x"04",x"8D",
    x"10",x"0F",x"79",x"0C",x"96",x"27",x"3B",x"BD",x"EB",x"7C",x"20",x"17",x"C6",x"49",x"8C",x"C6",
    x"4F",x"0D",x"8E",x"10",x"2B",x"40",x"33",x"86",x"10",x"C1",x"49",x"27",x"10",x"86",x"20",x"C1",
    x"4F",x"27",x"0A",x"C6",x"33",x"8C",x"C6",x"34",x"8C",x"C6",x"3C",x"0E",x"FB",x"97",x"90",x"D6",
    x"8E",x"BD",x"E3",x"A4",x"27",x"F3",x"AD",x"98",x"04",x"96",x"90",x"9A",x"8E",x"BD",x"E3",x"B0",
    x"A7",x"85",x"39",x"CC",x"02",x"00",x"20",x"3A",x"CC",x"00",x"FF",x"20",x"35",x"96",x"8E",x"81",
    x"02",x"26",x"04",x"0D",x"96",x"27",x"5B",x"0D",x"9A",x"26",x"03",x"BD",x"C4",x"24",x"7E",x"C3",
    x"81",x"DD",x"9C",x"DD",x"99",x"5C",x"D7",x"9B",x"BD",x"E0",x"F9",x"9D",x"B2",x"27",x"2A",x"9D",
    x"C2",x"81",x"2C",x"27",x"14",x"BD",x"CC",x"BA",x"9F",x"9C",x"20",x"0D",x"5F",x"80",x"4D",x"27",
    x"E0",x"4F",x"0F",x"9B",x"DD",x"99",x"BD",x"E0",x"76",x"9D",x"B2",x"27",x"0C",x"9D",x"C2",x"C6",
    x"52",x"9D",x"E0",x"26",x"AD",x"86",x"03",x"97",x"99",x"96",x"8E",x"2B",x"06",x"81",x"02",x"10",
    x"26",x"3F",x"A4",x"BD",x"E2",x"1C",x"DC",x"91",x"0D",x"9B",x"26",x"72",x"5D",x"26",x"9E",x"4D",
    x"27",x"03",x"7E",x"E2",x"33",x"0D",x"9A",x"26",x"F9",x"BD",x"C4",x"24",x"03",x"9E",x"8D",x"54",
    x"4C",x"97",x"7F",x"8D",x"48",x"D3",x"13",x"BD",x"C3",x"05",x"9E",x"13",x"BD",x"E3",x"62",x"D6",
    x"7A",x"26",x"04",x"A7",x"80",x"20",x"F5",x"9F",x"15",x"0D",x"7F",x"27",x"03",x"BD",x"E1",x"13",
    x"C6",x"03",x"6D",x"82",x"26",x"03",x"5A",x"26",x"F9",x"9E",x"15",x"9F",x"15",x"6F",x"80",x"5A",
    x"2A",x"F9",x"BD",x"E1",x"96",x"BD",x"C4",x"34",x"9E",x"13",x"BD",x"C3",x"FD",x"07",x"99",x"25",
    x"03",x"BD",x"E1",x"C6",x"07",x"99",x"10",x"25",x"FC",x"0C",x"7E",x"C3",x"7D",x"8D",x"00",x"8D",
    x"03",x"1E",x"89",x"39",x"8D",x"3C",x"0D",x"7A",x"27",x"F9",x"C6",x"35",x"0E",x"FB",x"5D",x"26",
    x"91",x"81",x"02",x"26",x"FA",x"8D",x"ED",x"34",x"02",x"8D",x"E2",x"1F",x"02",x"8D",x"DE",x"D3",
    x"9C",x"FD",x"22",x"3F",x"1F",x"01",x"A6",x"E0",x"27",x"0A",x"BD",x"E1",x"96",x"0D",x"99",x"27",
    x"D2",x"7E",x"E8",x"F6",x"8D",x"0C",x"D6",x"7A",x"26",x"D0",x"A7",x"80",x"31",x"3F",x"26",x"F4",
    x"20",x"D3",x"34",x"74",x"0F",x"7A",x"8D",x"43",x"10",x"2B",x"3E",x"F7",x"8D",x"34",x"AD",x"98",
    x"08",x"35",x"F4",x"34",x"76",x"8D",x"34",x"C5",x"10",x"27",x"04",x"C5",x"0F",x"26",x"0A",x"5D",
    x"10",x"2B",x"3E",x"DC",x"8D",x"1C",x"AD",x"98",x"0A",x"35",x"F6",x"34",x"16",x"0F",x"8F",x"8D",
    x"1A",x"10",x"2B",x"3E",x"D1",x"8D",x"0B",x"AD",x"98",x"0C",x"9F",x"7D",x"DD",x"7B",x"0D",x"7E",
    x"35",x"96",x"C4",x"0F",x"58",x"8E",x"23",x"C8",x"AE",x"85",x"39",x"8D",x"03",x"E6",x"85",x"39",
    x"8E",x"23",x"E8",x"D6",x"79",x"39",x"34",x"14",x"8D",x"F1",x"C4",x"8F",x"35",x"94",x"96",x"79",
    x"34",x"02",x"BD",x"E1",x"DA",x"8E",x"23",x"E8",x"6D",x"85",x"10",x"2B",x"3E",x"9B",x"8D",x"49",
    x"35",x"02",x"97",x"79",x"E6",x"85",x"8D",x"CA",x"AD",x"98",x"0E",x"7E",x"D5",x"DB",x"C6",x"24",
    x"9D",x"E0",x"BD",x"C7",x"2F",x"9D",x"E6",x"96",x"79",x"34",x"06",x"0F",x"79",x"9D",x"B2",x"81",
    x"29",x"27",x"03",x"BD",x"E1",x"CE",x"9D",x"DE",x"8D",x"1F",x"E6",x"61",x"BD",x"CB",x"ED",x"6C",
    x"61",x"6A",x"61",x"27",x"0A",x"BD",x"E3",x"62",x"BD",x"DD",x"02",x"A7",x"80",x"20",x"F2",x"35",
    x"06",x"97",x"79",x"7E",x"CB",x"85",x"86",x"20",x"8C",x"86",x"10",x"34",x"16",x"8D",x"91",x"27",
    x"0F",x"A6",x"85",x"27",x"0D",x"BD",x"22",x"87",x"84",x"30",x"A1",x"E4",x"10",x"26",x"FE",x"03",
    x"35",x"96",x"C6",x"39",x"0E",x"FB",x"9D",x"B2",x"5F",x"81",x"28",x"26",x"06",x"BD",x"C7",x"29",
    x"BD",x"CC",x"B2",x"96",x"79",x"34",x"02",x"5D",x"27",x"03",x"BD",x"E1",x"DD",x"8D",x"C7",x"9D",
    x"F3",x"35",x"02",x"97",x"79",x"D6",x"7D",x"0E",x"EC",x"00",x"16",x"28",x"29",x"2E",x"3A",x"FF",
    x"42",x"41",x"53",x"44",x"41",x"54",x"42",x"49",x"4E",x"F6",x"20",x"1B",x"0E",x"EC",x"0F",x"53",
    x"3F",x"0A",x"10",x"27",x"E7",x"0F",x"7E",x"CC",x"58",x"34",x"46",x"CE",x"A7",x"C1",x"CC",x"6E",
    x"6A",x"A7",x"C4",x"A6",x"C4",x"2A",x"0E",x"E7",x"C4",x"A6",x"C4",x"2B",x"16",x"86",x"64",x"A7",
    x"C4",x"A6",x"C4",x"2B",x"0E",x"3F",x"0A",x"27",x"FC",x"C1",x"02",x"27",x"F8",x"C1",x"03",x"10",
    x"27",x"E0",x"02",x"35",x"C6",x"AD",x"9F",x"22",x"55",x"8C",x"34",x"72",x"10",x"8E",x"24",x"45",
    x"E6",x"A4",x"27",x"09",x"A6",x"21",x"A7",x"A0",x"26",x"FA",x"5D",x"35",x"F2",x"3F",x"0A",x"2A",
    x"F9",x"CE",x"24",x"0E",x"A6",x"C5",x"2A",x"08",x"81",x"FF",x"27",x"D9",x"1F",x"89",x"1D",x"8C",
    x"8A",x"80",x"BD",x"DD",x"FD",x"20",x"D5",x"4B",x"59",x"42",x"44",x"E4",x"E7",x"E4",x"EB",x"E4",
    x"EC",x"E5",x"0A",x"E5",x"34",x"E4",x"F3",x"81",x"10",x"26",x"55",x"39",x"8D",x"BC",x"27",x"FC",
    x"1F",x"98",x"39",x"5F",x"39",x"53",x"43",x"52",x"4E",x"E5",x"05",x"E5",x"09",x"E4",x"EC",x"E5",
    x"0A",x"E5",x"34",x"E2",x"33",x"81",x"20",x"26",x"37",x"39",x"81",x"0D",x"26",x"09",x"7D",x"20",
    x"2C",x"27",x"04",x"C6",x"18",x"8D",x"1B",x"F6",x"20",x"2A",x"54",x"24",x"13",x"34",x"02",x"B6",
    x"20",x"1B",x"4A",x"2B",x"03",x"BD",x"ED",x"B8",x"35",x"02",x"81",x"0A",x"26",x"02",x"8D",x"00",
    x"1F",x"89",x"3F",x"82",x"B6",x"20",x"1C",x"4A",x"C6",x"28",x"1F",x"01",x"CC",x"0D",x"1A",x"39",
    x"7E",x"E2",x"33",x"4C",x"50",x"52",x"54",x"E5",x"53",x"E5",x"83",x"E2",x"33",x"E5",x"70",x"E5",
    x"A8",x"E2",x"33",x"8D",x"B0",x"0D",x"8C",x"10",x"26",x"06",x"37",x"CE",x"24",x"06",x"8D",x"4F",
    x"03",x"8C",x"C6",x"04",x"F7",x"20",x"42",x"3F",x"24",x"24",x"0F",x"8D",x"18",x"7E",x"EB",x"8F",
    x"0D",x"AB",x"26",x"04",x"81",x"16",x"26",x"03",x"03",x"AB",x"39",x"81",x"0D",x"26",x"0C",x"0F",
    x"89",x"20",x"1C",x"8D",x"54",x"0F",x"8C",x"C6",x"10",x"20",x"D9",x"81",x"20",x"25",x"10",x"D6",
    x"89",x"D1",x"8A",x"25",x"08",x"34",x"02",x"8D",x"44",x"35",x"02",x"0F",x"89",x"0C",x"89",x"C6",
    x"01",x"F7",x"20",x"42",x"1F",x"89",x"20",x"BF",x"9E",x"89",x"86",x"0D",x"D6",x"8B",x"39",x"0F",
    x"89",x"C6",x"28",x"A6",x"C4",x"27",x"14",x"9E",x"B3",x"34",x"10",x"DF",x"B3",x"9D",x"B2",x"BD",
    x"C6",x"4B",x"DC",x"28",x"4D",x"26",x"53",x"35",x"10",x"9F",x"B3",x"D7",x"8A",x"4F",x"8B",x"0D",
    x"91",x"8A",x"23",x"FA",x"80",x"1A",x"97",x"8B",x"39",x"0D",x"89",x"27",x"9D",x"0F",x"89",x"86",
    x"0D",x"8D",x"BC",x"86",x"0A",x"20",x"B8",x"9D",x"AC",x"96",x"8C",x"34",x"02",x"26",x"03",x"17",
    x"FF",x"6E",x"8D",x"E5",x"C6",x"02",x"17",x"FF",x"6B",x"A6",x"E0",x"27",x"86",x"39",x"BD",x"E7",
    x"75",x"BD",x"ED",x"D0",x"9D",x"B2",x"27",x"F5",x"8D",x"08",x"10",x"27",x"07",x"B7",x"C6",x"14",
    x"3F",x"82",x"9D",x"C2",x"9D",x"E6",x"C1",x"01",x"23",x"E3",x"0E",x"F6",x"C6",x"02",x"8D",x"02",
    x"C6",x"01",x"BD",x"E6",x"A4",x"27",x"15",x"34",x"04",x"53",x"F4",x"20",x"2A",x"34",x"04",x"8D",
    x"E3",x"27",x"02",x"6F",x"61",x"35",x"04",x"EA",x"E0",x"F7",x"20",x"2A",x"BD",x"E7",x"04",x"39",
    x"F6",x"20",x"1E",x"81",x"2C",x"27",x"06",x"9D",x"E6",x"C1",x"18",x"22",x"CD",x"34",x"04",x"F6",
    x"20",x"20",x"9D",x"B2",x"27",x"0F",x"9D",x"C2",x"F6",x"20",x"20",x"81",x"2C",x"27",x"06",x"9D",
    x"E6",x"C1",x"18",x"22",x"B5",x"E1",x"E4",x"25",x"B1",x"8D",x"1E",x"35",x"04",x"8D",x"17",x"8D",
    x"CB",x"27",x"06",x"8D",x"9F",x"CB",x"74",x"8D",x"0B",x"8D",x"29",x"BD",x"CC",x"AB",x"C1",x"02",
    x"22",x"C9",x"CB",x"78",x"20",x"6A",x"86",x"20",x"8C",x"86",x"10",x"34",x"02",x"86",x"FF",x"4C",
    x"C0",x"0A",x"24",x"FB",x"CB",x"0A",x"AA",x"E4",x"EA",x"E0",x"34",x"06",x"C6",x"1F",x"8D",x"62",
    x"35",x"04",x"20",x"5A",x"9D",x"B2",x"26",x"62",x"35",x"86",x"9D",x"AC",x"81",x"AB",x"10",x"27",
    x"FF",x"35",x"C6",x"5F",x"D7",x"9F",x"8D",x"EC",x"27",x"06",x"8D",x"51",x"CA",x"40",x"8D",x"32",
    x"8D",x"42",x"27",x"06",x"8D",x"47",x"CA",x"50",x"8D",x"28",x"0D",x"9F",x"27",x"0C",x"8D",x"34",
    x"27",x"08",x"8D",x"39",x"CA",x"60",x"8D",x"18",x"03",x"9F",x"8D",x"28",x"27",x"07",x"BD",x"E6",
    x"14",x"C6",x"7B",x"8D",x"0D",x"0D",x"9F",x"27",x"2A",x"8D",x"B9",x"BD",x"E6",x"12",x"CB",x"76",
    x"0F",x"9F",x"34",x"04",x"C6",x"1B",x"8D",x"0A",x"0D",x"9F",x"27",x"04",x"C6",x"20",x"8D",x"02",
    x"35",x"04",x"3F",x"82",x"9D",x"B2",x"27",x"A0",x"9D",x"C2",x"81",x"2C",x"39",x"9D",x"E6",x"C1",
    x"0F",x"22",x"36",x"39",x"8D",x"58",x"3F",x"14",x"7E",x"D5",x"DB",x"8D",x"51",x"8D",x"58",x"3F",
    x"1A",x"C1",x"16",x"26",x"22",x"3F",x"1A",x"86",x"7B",x"CE",x"F6",x"4D",x"4C",x"33",x"43",x"E1",
    x"C4",x"26",x"F9",x"3F",x"1A",x"CE",x"EA",x"AD",x"8B",x"04",x"81",x"80",x"27",x"04",x"E1",x"C0",
    x"22",x"F6",x"1F",x"89",x"27",x"01",x"5F",x"0E",x"EC",x"0E",x"F6",x"CC",x"01",x"3F",x"8D",x"0D",
    x"34",x"06",x"9D",x"C2",x"CC",x"00",x"C7",x"8D",x"04",x"1F",x"02",x"35",x"90",x"DD",x"67",x"BD",
    x"C9",x"85",x"10",x"93",x"67",x"23",x"02",x"DC",x"67",x"39",x"C6",x"C8",x"9D",x"E0",x"BD",x"C7",
    x"2F",x"8D",x"D8",x"0E",x"DE",x"8D",x"D4",x"30",x"01",x"8C",x"00",x"28",x"23",x"03",x"8E",x"00",
    x"28",x"10",x"8C",x"00",x"18",x"23",x"04",x"10",x"8E",x"00",x"18",x"1F",x"20",x"34",x"04",x"1F",
    x"10",x"35",x"82",x"8D",x"D9",x"8D",x"32",x"39",x"9D",x"C2",x"9D",x"CD",x"BD",x"D6",x"27",x"10",
    x"83",x"FF",x"F0",x"2D",x"A4",x"10",x"83",x"00",x"0F",x"2E",x"9E",x"20",x"64",x"37",x"30",x"8D",
    x"C6",x"36",x"30",x"39",x"CE",x"25",x"81",x"37",x"30",x"81",x"C8",x"27",x"02",x"8D",x"AF",x"CE",
    x"25",x"81",x"36",x"30",x"34",x"30",x"8D",x"A2",x"8C",x"34",x"30",x"CE",x"25",x"85",x"36",x"30",
    x"9D",x"B2",x"27",x"36",x"81",x"2C",x"27",x"C0",x"BD",x"CC",x"15",x"F7",x"20",x"36",x"9D",x"B2",
    x"27",x"05",x"9D",x"C2",x"BD",x"E6",x"B3",x"CE",x"25",x"7D",x"8D",x"C1",x"33",x"44",x"8D",x"BD",
    x"35",x"70",x"B6",x"20",x"2A",x"34",x"02",x"84",x"FC",x"8D",x"07",x"BD",x"E7",x"77",x"8D",x"06",
    x"35",x"02",x"B7",x"20",x"2A",x"39",x"34",x"40",x"3F",x"92",x"F6",x"20",x"2B",x"54",x"54",x"54",
    x"54",x"F7",x"20",x"29",x"35",x"30",x"7F",x"20",x"36",x"3F",x"90",x"81",x"FF",x"10",x"27",x"F4",
    x"60",x"8D",x"91",x"BE",x"25",x"81",x"10",x"BE",x"25",x"83",x"3F",x"8E",x"0F",x"A0",x"81",x"46",
    x"26",x"04",x"97",x"A0",x"9D",x"AC",x"BD",x"E7",x"B4",x"CE",x"25",x"7D",x"96",x"A0",x"26",x"0F",
    x"AE",x"44",x"8D",x"E6",x"8D",x"E0",x"AE",x"C4",x"8D",x"E0",x"10",x"AE",x"42",x"20",x"DB",x"10",
    x"AE",x"42",x"AE",x"C4",x"8D",x"C3",x"AE",x"44",x"8D",x"D0",x"10",x"AC",x"46",x"27",x"A6",x"22",
    x"03",x"31",x"21",x"8C",x"31",x"3F",x"20",x"EA",x"BD",x"22",x"75",x"C6",x"FF",x"9D",x"E0",x"C6",
    x"99",x"9D",x"E0",x"BD",x"C7",x"29",x"C6",x"D4",x"9D",x"E0",x"BD",x"CC",x"B2",x"D1",x"AA",x"24",
    x"1C",x"86",x"08",x"3D",x"D3",x"1F",x"1F",x"01",x"30",x"09",x"86",x"08",x"34",x"12",x"9D",x"E6",
    x"35",x"12",x"E7",x"82",x"4A",x"27",x"51",x"34",x"12",x"9D",x"C2",x"20",x"F1",x"0E",x"F6",x"8D",
    x"02",x"0E",x"EC",x"BD",x"CC",x"B2",x"BD",x"E6",x"16",x"1F",x"98",x"3F",x"9C",x"3F",x"16",x"20",
    x"02",x"8D",x"F0",x"C6",x"00",x"C2",x"00",x"7E",x"D5",x"DB",x"9D",x"AC",x"BD",x"E4",x"79",x"3F",
    x"16",x"24",x"F9",x"8D",x"1A",x"34",x"30",x"9D",x"F0",x"35",x"06",x"8D",x"06",x"9D",x"C2",x"9D",
    x"F0",x"35",x"06",x"9D",x"ED",x"96",x"39",x"BD",x"D6",x"65",x"9E",x"37",x"7E",x"D7",x"F3",x"3F",
    x"18",x"24",x"05",x"8E",x"FF",x"FF",x"1F",x"12",x"39",x"BD",x"E1",x"01",x"9D",x"B2",x"27",x"06",
    x"BD",x"CC",x"BA",x"BF",x"22",x"3F",x"6E",x"9F",x"22",x"3F",x"3F",x"88",x"C6",x"0C",x"3F",x"82",
    x"8D",x"FA",x"3F",x"0A",x"3F",x"16",x"24",x"18",x"3F",x"18",x"25",x"14",x"9F",x"32",x"10",x"8E",
    x"00",x"C8",x"3F",x"0E",x"C1",x"08",x"26",x"02",x"0C",x"78",x"C1",x"09",x"26",x"02",x"0A",x"78",
    x"03",x"29",x"10",x"8E",x"00",x"00",x"3F",x"0E",x"03",x"29",x"C1",x"0D",x"26",x"D4",x"35",x"04",
    x"D7",x"19",x"35",x"88",x"12",x"C6",x"21",x"1F",x"9B",x"0F",x"05",x"C6",x"1B",x"3F",x"02",x"CC",
    x"46",x"66",x"B7",x"20",x"2B",x"3F",x"02",x"8D",x"B3",x"C6",x"A5",x"F1",x"22",x"00",x"27",x"1E",
    x"8E",x"E9",x"35",x"BF",x"00",x"1E",x"7D",x"20",x"80",x"27",x"02",x"3F",x"A8",x"10",x"CE",x"5F",
    x"FF",x"8D",x"26",x"8E",x"EA",x"89",x"BD",x"CE",x"2C",x"BD",x"C4",x"24",x"20",x"13",x"10",x"DE",
    x"19",x"D6",x"9E",x"27",x"03",x"BD",x"C4",x"24",x"BD",x"C4",x"39",x"BD",x"E1",x"C6",x"BD",x"22",
    x"8A",x"1C",x"AF",x"BD",x"ED",x"C5",x"7E",x"C3",x"7D",x"8E",x"21",x"00",x"6F",x"80",x"8C",x"25",
    x"A3",x"23",x"F9",x"9F",x"13",x"F7",x"22",x"00",x"8C",x"63",x"80",x"A6",x"84",x"43",x"A7",x"84",
    x"A1",x"84",x"27",x"F5",x"30",x"1E",x"9F",x"A1",x"9F",x"1F",x"9F",x"1B",x"30",x"89",x"FE",x"D4",
    x"9F",x"19",x"86",x"02",x"97",x"8D",x"8E",x"EA",x"2C",x"CE",x"22",x"01",x"C6",x"0A",x"8D",x"5A",
    x"8E",x"21",x"F9",x"AF",x"43",x"AF",x"48",x"CE",x"22",x"33",x"CC",x"7E",x"04",x"8D",x"31",x"8E",
    x"21",x"F6",x"C6",x"0C",x"AF",x"C1",x"5A",x"26",x"FB",x"C6",x"01",x"8D",x"23",x"8E",x"E2",x"39",
    x"C6",x"07",x"8D",x"1C",x"CC",x"39",x"0B",x"8D",x"17",x"8E",x"EA",x"BA",x"CE",x"23",x"90",x"C6",
    x"40",x"8D",x"27",x"73",x"24",x"4E",x"8E",x"EA",x"36",x"CE",x"21",x"AC",x"C6",x"54",x"20",x"1A",
    x"A7",x"C0",x"AF",x"C1",x"5A",x"26",x"F9",x"39",x"8D",x"18",x"6F",x"01",x"30",x"1F",x"9C",x"1F",
    x"24",x"F8",x"8E",x"EA",x"B3",x"CE",x"20",x"39",x"C6",x"07",x"A6",x"80",x"A7",x"C0",x"5A",x"26",
    x"F9",x"39",x"9E",x"1F",x"D6",x"AA",x"86",x"08",x"3D",x"30",x"8B",x"39",x"56",x"C0",x"A0",x"C2",
    x"5F",x"27",x"C1",x"CC",x"C0",x"00",x"0C",x"B4",x"26",x"02",x"0C",x"B3",x"B6",x"00",x"00",x"81",
    x"20",x"27",x"F3",x"81",x"3A",x"24",x"04",x"80",x"30",x"80",x"D0",x"39",x"7E",x"C7",x"32",x"96",
    x"4B",x"7E",x"D8",x"21",x"7E",x"D8",x"29",x"9D",x"CA",x"9D",x"DB",x"7E",x"D6",x"58",x"9D",x"DB",
    x"7E",x"D6",x"60",x"9D",x"CA",x"7E",x"C7",x"42",x"C6",x"29",x"7E",x"C7",x"34",x"7E",x"E3",x"73",
    x"7E",x"CC",x"B0",x"7E",x"D6",x"6B",x"4F",x"7E",x"D5",x"DC",x"7E",x"C8",x"AA",x"7E",x"E3",x"8B",
    x"C6",x"05",x"8C",x"C6",x"02",x"7E",x"C3",x"24",x"00",x"00",x"0C",x"4D",x"4F",x"20",x"42",x"41",
    x"53",x"49",x"43",x"20",x"31",x"2E",x"30",x"20",x"0A",x"0D",x"28",x"63",x"29",x"20",x"4D",x"69",
    x"63",x"72",x"6F",x"73",x"6F",x"66",x"74",x"20",x"31",x"39",x"38",x"34",x"00",x"61",x"65",x"69",
    x"6F",x"75",x"FF",x"00",x"05",x"00",x"18",x"00",x"00",x"02",x"9D",x"2E",x"06",x"A2",x"1D",x"1E",
    x"2C",x"83",x"99",x"A0",x"28",x"34",x"0B",x"25",x"10",x"22",x"9A",x"0A",x"1C",x"2A",x"A4",x"26",
    x"21",x"03",x"9C",x"05",x"0F",x"1F",x"1B",x"20",x"11",x"24",x"9B",x"98",x"08",x"16",x"01",x"2D",
    x"39",x"8A",x"A1",x"97",x"3B",x"09",x"07",x"9F",x"33",x"2B",x"37",x"A6",x"46",x"04",x"3C",x"44",
    x"32",x"02",x"E4",x"D7",x"E4",x"F5",x"EA",x"FA",x"E5",x"43",x"43",x"41",x"53",x"53",x"EB",x"31",
    x"EB",x"6A",x"EB",x"2A",x"EB",x"9E",x"EB",x"0A",x"EB",x"22",x"03",x"8F",x"CC",x"01",x"00",x"9E",
    x"FE",x"39",x"D6",x"94",x"E0",x"3F",x"A6",x"AB",x"6A",x"3F",x"26",x"14",x"34",x"02",x"8D",x"62",
    x"35",x"82",x"8D",x"72",x"26",x"01",x"43",x"1E",x"89",x"39",x"8D",x"6A",x"26",x"E4",x"03",x"7A",
    x"39",x"0D",x"95",x"26",x"5D",x"81",x"10",x"27",x"7B",x"8E",x"23",x"FA",x"6D",x"80",x"10",x"27",
    x"F4",x"DE",x"CE",x"22",x"91",x"C6",x"0B",x"BD",x"EA",x"1A",x"DC",x"91",x"ED",x"C1",x"96",x"96",
    x"A7",x"C0",x"C6",x"0E",x"E7",x"51",x"86",x"02",x"97",x"95",x"0F",x"93",x"D7",x"97",x"BD",x"EC",
    x"00",x"96",x"96",x"97",x"97",x"8D",x"2F",x"6F",x"3F",x"39",x"0D",x"95",x"27",x"13",x"81",x"20",
    x"26",x"0A",x"8D",x"22",x"27",x"02",x"8D",x"4E",x"C6",x"FF",x"8D",x"4C",x"BD",x"EC",x"1E",x"0F",
    x"95",x"39",x"8D",x"64",x"27",x"07",x"2B",x"04",x"8D",x"0C",x"27",x"F6",x"39",x"8D",x"ED",x"C6",
    x"35",x"8C",x"C6",x"3B",x"0E",x"FB",x"10",x"8E",x"22",x"91",x"4F",x"E6",x"3F",x"39",x"34",x"02",
    x"8D",x"F4",x"CB",x"02",x"26",x"04",x"8D",x"1E",x"C6",x"02",x"5A",x"E7",x"3F",x"31",x"AB",x"35",
    x"02",x"A7",x"3F",x"39",x"8D",x"7C",x"8D",x"AD",x"EC",x"2B",x"DD",x"91",x"A6",x"2D",x"97",x"96",
    x"97",x"97",x"0C",x"95",x"20",x"BC",x"C6",x"01",x"D7",x"93",x"8D",x"34",x"20",x"97",x"86",x"02",
    x"CE",x"E4",x"60",x"BD",x"DF",x"96",x"96",x"8E",x"81",x"02",x"10",x"26",x"36",x"18",x"8D",x"D4",
    x"0D",x"93",x"2B",x"98",x"8D",x"9C",x"20",x"F8",x"8D",x"3F",x"10",x"8E",x"22",x"90",x"3F",x"20",
    x"4D",x"26",x"9A",x"A6",x"A0",x"80",x"02",x"97",x"94",x"A7",x"3F",x"8D",x"1D",x"D7",x"93",x"39",
    x"8D",x"27",x"8D",x"92",x"30",x"A4",x"5D",x"27",x"05",x"AB",x"80",x"5A",x"26",x"FB",x"40",x"A7",
    x"84",x"6C",x"A2",x"6C",x"A4",x"4F",x"D6",x"93",x"3F",x"20",x"0D",x"97",x"27",x"13",x"4F",x"97",
    x"05",x"3F",x"22",x"24",x"0C",x"C6",x"3C",x"0E",x"FB",x"96",x"95",x"8A",x"01",x"0D",x"05",x"27",
    x"EE",x"39",x"96",x"24",x"4C",x"97",x"98",x"8E",x"EC",x"8E",x"8D",x"22",x"0F",x"97",x"8D",x"A8",
    x"26",x"FA",x"8D",x"DA",x"8E",x"23",x"FA",x"6D",x"80",x"27",x"0B",x"C6",x"0B",x"A6",x"80",x"A1",
    x"A0",x"26",x"12",x"5A",x"26",x"F7",x"8E",x"EC",x"9C",x"8D",x"1F",x"8E",x"EC",x"99",x"0D",x"98",
    x"26",x"CF",x"7E",x"CE",x"2C",x"8E",x"EC",x"A4",x"8D",x"10",x"20",x"CB",x"1F",x"89",x"9D",x"AC",
    x"C1",x"96",x"27",x"B5",x"C1",x"C3",x"27",x"A6",x"0E",x"F9",x"8D",x"E2",x"0D",x"98",x"26",x"E0",
    x"8E",x"22",x"91",x"C6",x"08",x"8D",x"05",x"BD",x"CE",x"3E",x"C6",x"03",x"7E",x"CE",x"32",x"0D",
    x"0A",x"53",x"65",x"61",x"72",x"63",x"68",x"69",x"6E",x"67",x"0D",x"0A",x"00",x"46",x"6F",x"75",
    x"6E",x"64",x"3A",x"20",x"00",x"53",x"6B",x"69",x"70",x"3A",x"20",x"00",x"8E",x"24",x"52",x"BD",
    x"E3",x"62",x"0D",x"7A",x"26",x"13",x"81",x"0D",x"27",x"0F",x"81",x"16",x"27",x"04",x"81",x"20",
    x"25",x"ED",x"A7",x"80",x"8C",x"25",x"51",x"25",x"E6",x"BD",x"22",x"7E",x"7E",x"ED",x"7A",x"BD",
    x"E3",x"B6",x"26",x"D8",x"C6",x"70",x"BD",x"E6",x"F0",x"B6",x"20",x"1E",x"F6",x"20",x"20",x"DD",
    x"84",x"8D",x"3A",x"DD",x"82",x"8D",x"76",x"96",x"84",x"8D",x"72",x"96",x"85",x"8D",x"6E",x"BD",
    x"ED",x"C5",x"8D",x"73",x"BD",x"E6",x"0E",x"81",x"03",x"27",x"72",x"81",x"0D",x"27",x"22",x"BD",
    x"EE",x"3F",x"C6",x"0B",x"8E",x"EF",x"01",x"EE",x"81",x"A1",x"80",x"27",x"0A",x"5A",x"26",x"F7",
    x"81",x"20",x"25",x"DB",x"CE",x"ED",x"98",x"8D",x"04",x"AD",x"C4",x"20",x"D2",x"FC",x"20",x"1B",
    x"39",x"BD",x"EE",x"45",x"91",x"82",x"26",x"02",x"DC",x"82",x"34",x"06",x"BD",x"EE",x"61",x"DD",
    x"80",x"EC",x"E4",x"8E",x"24",x"52",x"10",x"93",x"80",x"22",x"39",x"BD",x"EE",x"DE",x"8C",x"25",
    x"51",x"27",x"31",x"C1",x"16",x"26",x"0B",x"8C",x"25",x"4E",x"27",x"28",x"E7",x"80",x"DC",x"87",
    x"A7",x"80",x"E7",x"80",x"EC",x"E4",x"BD",x"EE",x"51",x"ED",x"E4",x"20",x"D9",x"4A",x"2B",x"04",
    x"8D",x"56",x"63",x"86",x"39",x"8D",x"45",x"BD",x"E3",x"62",x"97",x"86",x"39",x"8D",x"50",x"BD",
    x"CD",x"F0",x"43",x"39",x"AF",x"E4",x"8D",x"F5",x"35",x"10",x"6F",x"80",x"8E",x"24",x"51",x"39",
    x"5A",x"26",x"29",x"91",x"84",x"26",x"25",x"39",x"8D",x"42",x"C1",x"28",x"26",x"1E",x"91",x"85",
    x"20",x"F3",x"8D",x"D1",x"8D",x"CF",x"8D",x"85",x"91",x"82",x"26",x"06",x"D1",x"83",x"24",x"02",
    x"D7",x"83",x"C1",x"28",x"26",x"06",x"8D",x"6B",x"27",x"02",x"8D",x"36",x"D6",x"86",x"3F",x"02",
    x"34",x"12",x"96",x"85",x"8D",x"AA",x"35",x"92",x"8E",x"20",x"00",x"6F",x"86",x"39",x"12",x"8D",
    x"7F",x"8D",x"46",x"8D",x"0B",x"C6",x"11",x"8C",x"CA",x"40",x"3F",x"82",x"96",x"84",x"C6",x"01",
    x"DD",x"80",x"34",x"06",x"C6",x"1F",x"3F",x"02",x"D6",x"80",x"8D",x"EC",x"D6",x"81",x"8D",x"E8",
    x"35",x"86",x"34",x"06",x"8D",x"7B",x"91",x"85",x"22",x"51",x"DD",x"80",x"8D",x"57",x"D6",x"80",
    x"91",x"84",x"25",x"47",x"27",x"23",x"91",x"82",x"26",x"02",x"0A",x"82",x"6A",x"E4",x"33",x"C9",
    x"FF",x"00",x"BD",x"E6",x"89",x"86",x"0A",x"20",x"1C",x"FC",x"20",x"1B",x"4A",x"4C",x"8D",x"03",
    x"27",x"FB",x"39",x"8E",x"20",x"00",x"6D",x"86",x"39",x"D1",x"85",x"24",x"1E",x"5C",x"D7",x"80",
    x"BD",x"E6",x"86",x"86",x"0B",x"8D",x"19",x"1F",x"89",x"8D",x"4C",x"B6",x"20",x"1B",x"4A",x"8D",
    x"87",x"D6",x"84",x"BD",x"E6",x"86",x"D6",x"85",x"BD",x"E6",x"89",x"35",x"06",x"8D",x"91",x"C6",
    x"5F",x"F7",x"20",x"2C",x"39",x"FC",x"20",x"1B",x"4A",x"2B",x"04",x"8D",x"C6",x"27",x"F9",x"4C",
    x"5F",x"5C",x"C1",x"29",x"27",x"F9",x"39",x"4A",x"91",x"84",x"2D",x"F3",x"8D",x"B5",x"26",x"EF",
    x"8C",x"8D",x"A6",x"C6",x"29",x"5A",x"27",x"EF",x"34",x"06",x"8D",x"72",x"C1",x"20",x"35",x"06",
    x"27",x"F3",x"39",x"32",x"62",x"C6",x"20",x"8D",x"03",x"BD",x"ED",x"AE",x"7E",x"ED",x"D2",x"34",
    x"06",x"8D",x"DE",x"10",x"A3",x"E4",x"25",x"E6",x"91",x"85",x"26",x"05",x"C1",x"28",x"26",x"01",
    x"5A",x"8D",x"80",x"27",x"11",x"C1",x"27",x"26",x"0D",x"1F",x"03",x"35",x"06",x"BD",x"ED",x"E2",
    x"DC",x"80",x"34",x"06",x"1F",x"30",x"10",x"A3",x"E4",x"2B",x"C8",x"DD",x"80",x"C6",x"09",x"8D",
    x"46",x"DC",x"80",x"5A",x"26",x"F0",x"C6",x"28",x"4A",x"20",x"EB",x"34",x"06",x"DD",x"80",x"8D",
    x"A0",x"1F",x"01",x"9C",x"80",x"25",x"2E",x"9C",x"80",x"23",x"0C",x"DC",x"80",x"8D",x"82",x"DD",
    x"80",x"C6",x"08",x"8D",x"22",x"20",x"F0",x"8D",x"9C",x"35",x"06",x"7E",x"ED",x"D0",x"34",x"10",
    x"1F",x"01",x"4F",x"1E",x"01",x"3F",x"1A",x"C1",x"16",x"26",x"0A",x"3F",x"1A",x"D7",x"87",x"3F",
    x"1A",x"D7",x"88",x"C6",x"16",x"35",x"90",x"8D",x"83",x"CE",x"FF",x"FF",x"FF",x"20",x"2E",x"3F",
    x"82",x"ED",x"83",x"0B",x"ED",x"8E",x"0A",x"ED",x"8A",x"09",x"ED",x"80",x"08",x"ED",x"AC",x"18",
    x"ED",x"92",x"16",x"ED",x"88",x"0C",x"EE",x"7F",x"1C",x"EE",x"BB",x"1D",x"ED",x"CC",x"1E",x"ED",
    x"B8",x"17",x"9D",x"B2",x"27",x"76",x"9D",x"C2",x"BD",x"CB",x"F5",x"31",x"84",x"D7",x"02",x"0D",
    x"02",x"27",x"EF",x"8D",x"68",x"81",x"20",x"27",x"F6",x"81",x"3B",x"27",x"F2",x"8D",x"02",x"20",
    x"EE",x"5F",x"81",x"50",x"27",x"6F",x"8E",x"EF",x"DB",x"0D",x"02",x"27",x"0E",x"E6",x"A4",x"30",
    x"12",x"10",x"A3",x"81",x"27",x"51",x"8C",x"EF",x"DB",x"26",x"F6",x"A1",x"84",x"27",x"09",x"30",
    x"05",x"8C",x"EF",x"CD",x"26",x"F5",x"0E",x"F6",x"8D",x"33",x"24",x"FA",x"5F",x"80",x"30",x"34",
    x"02",x"86",x"0A",x"3D",x"4D",x"26",x"EF",x"EB",x"E0",x"25",x"EB",x"0D",x"02",x"27",x"08",x"8D",
    x"1C",x"25",x"EA",x"31",x"3F",x"0C",x"02",x"E1",x"01",x"25",x"DB",x"E1",x"02",x"22",x"D7",x"8C",
    x"EF",x"EA",x"26",x"05",x"CE",x"FF",x"41",x"E6",x"C5",x"E7",x"98",x"03",x"39",x"0D",x"02",x"27",
    x"C5",x"A6",x"A0",x"0A",x"02",x"0E",x"B9",x"8D",x"F4",x"1F",x"10",x"83",x"EF",x"CE",x"C1",x"05",
    x"23",x"01",x"5A",x"0D",x"02",x"27",x"14",x"A6",x"A4",x"81",x"23",x"26",x"03",x"5C",x"8D",x"DD",
    x"81",x"62",x"26",x"07",x"8D",x"D7",x"5A",x"26",x"02",x"C6",x"0C",x"3F",x"9E",x"44",x"4F",x"52",
    x"45",x"4D",x"49",x"46",x"41",x"53",x"4F",x"4C",x"41",x"53",x"49",x"54",x"01",x"FF",x"20",x"3A",
    x"41",x"00",x"FF",x"20",x"3D",x"4C",x"01",x"60",x"20",x"3C",x"4F",x"01",x"05",x"20",x"3F",x"9C",
    x"19",x"25",x"03",x"11",x"93",x"15",x"10",x"25",x"32",x"8A",x"7E",x"FF",x"E4",x"FD",x"E9",x"35");

  CONSTANT ROM_BASIC6_1 : arr8 := (
    x"3F",x"04",x"86",x"A5",x"B1",x"1F",x"DF",x"27",x"45",x"B7",x"1F",x"DF",x"86",x"0F",x"CE",x"1F",
    x"E0",x"10",x"8E",x"00",x"00",x"8E",x"1F",x"FF",x"3F",x"3C",x"48",x"AF",x"C6",x"8E",x"10",x"00",
    x"CE",x"C0",x"2E",x"10",x"AE",x"C6",x"44",x"3F",x"3C",x"4A",x"2A",x"E2",x"20",x"20",x"00",x"00",
    x"00",x"00",x"00",x"00",x"03",x"AA",x"04",x"20",x"00",x"00",x"0F",x"F0",x"0F",x"FF",x"0E",x"E7",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"8E",x"C4",
    x"5E",x"9F",x"70",x"8E",x"C2",x"3C",x"BD",x"FB",x"FE",x"BD",x"C1",x"2C",x"BD",x"FB",x"99",x"43",
    x"26",x"04",x"5F",x"7E",x"C1",x"1B",x"8E",x"C3",x"05",x"C6",x"01",x"BD",x"FB",x"F8",x"B6",x"A0",
    x"00",x"81",x"52",x"26",x"03",x"8E",x"C3",x"35",x"C6",x"02",x"BD",x"FB",x"F8",x"8E",x"C3",x"40",
    x"C6",x"03",x"BD",x"FB",x"F8",x"86",x"04",x"B7",x"A7",x"E5",x"CC",x"55",x"13",x"8E",x"6F",x"E0",
    x"AB",x"85",x"5A",x"2A",x"FB",x"B1",x"6F",x"F5",x"26",x"11",x"C6",x"04",x"BD",x"FB",x"F8",x"8E",
    x"C3",x"5C",x"BD",x"FB",x"FE",x"86",x"80",x"9A",x"7F",x"97",x"7F",x"86",x"02",x"B7",x"A7",x"E5",
    x"8E",x"C3",x"5F",x"BD",x"FB",x"FE",x"86",x"24",x"8D",x"74",x"96",x"79",x"85",x"C0",x"26",x"03",
    x"BD",x"CE",x"A6",x"C6",x"34",x"F7",x"A7",x"C1",x"F6",x"A7",x"C1",x"2B",x"16",x"C6",x"28",x"F7",
    x"A7",x"C1",x"F6",x"A7",x"C1",x"2B",x"0C",x"C6",x"0E",x"F7",x"A7",x"C1",x"F6",x"A7",x"C1",x"10",
    x"2A",x"0E",x"18",x"3F",x"0A",x"5D",x"27",x"04",x"C0",x"30",x"20",x"16",x"BD",x"C1",x"72",x"25",
    x"C9",x"3F",x"16",x"24",x"C5",x"81",x"04",x"24",x"C1",x"C0",x"10",x"04",x"7F",x"25",x"01",x"5C",
    x"09",x"7F",x"C1",x"04",x"22",x"B4",x"26",x"04",x"0D",x"7F",x"2A",x"AE",x"C1",x"03",x"27",x"26",
    x"5D",x"26",x"08",x"04",x"7F",x"25",x"04",x"09",x"7F",x"20",x"9F",x"8D",x"03",x"7E",x"F1",x"97",
    x"3F",x"04",x"7F",x"1F",x"DF",x"8E",x"1F",x"E0",x"86",x"FF",x"3F",x"BC",x"86",x"28",x"C6",x"60",
    x"3F",x"02",x"4A",x"26",x"FB",x"39",x"17",x"00",x"BF",x"3F",x"0A",x"C0",x"31",x"C1",x"03",x"23",
    x"12",x"8D",x"30",x"25",x"F4",x"3F",x"16",x"24",x"F0",x"81",x"04",x"24",x"EC",x"C0",x"10",x"C1",
    x"03",x"22",x"E6",x"CE",x"C1",x"5B",x"58",x"AD",x"D5",x"20",x"DB",x"C8",x"98",x"C1",x"68",x"C1",
    x"6B",x"C1",x"63",x"32",x"62",x"7E",x"C0",x"4E",x"C6",x"04",x"8C",x"C6",x"80",x"D8",x"79",x"D7",
    x"79",x"39",x"86",x"4F",x"3F",x"18",x"25",x"F9",x"4D",x"26",x"05",x"17",x"00",x"3A",x"25",x"F1",
    x"1F",x"20",x"54",x"54",x"54",x"34",x"06",x"58",x"86",x"A0",x"3D",x"34",x"06",x"1F",x"10",x"44",
    x"56",x"54",x"54",x"E7",x"62",x"E3",x"E1",x"1F",x"02",x"8D",x"0B",x"8E",x"09",x"C4",x"BD",x"F4",
    x"75",x"8D",x"03",x"4F",x"35",x"86",x"34",x"20",x"3F",x"06",x"86",x"08",x"63",x"A4",x"31",x"A8",
    x"28",x"4A",x"26",x"F8",x"35",x"A0",x"4F",x"39",x"10",x"8C",x"00",x"28",x"23",x"F8",x"10",x"8C",
    x"00",x"58",x"24",x"F2",x"3F",x"16",x"24",x"EE",x"9F",x"32",x"10",x"8E",x"00",x"28",x"10",x"9F",
    x"34",x"10",x"8E",x"00",x"57",x"0F",x"29",x"3F",x"0E",x"3F",x"0A",x"C1",x"08",x"26",x"02",x"0C",
    x"78",x"C1",x"09",x"26",x"02",x"0A",x"78",x"C6",x"F9",x"D7",x"29",x"0C",x"35",x"10",x"8E",x"00",
    x"28",x"3F",x"0E",x"3F",x"18",x"24",x"C1",x"39",x"8E",x"C3",x"66",x"BD",x"FB",x"FE",x"17",x"FF",
    x"2B",x"C6",x"01",x"8E",x"C3",x"B0",x"BD",x"FB",x"F8",x"C6",x"02",x"8E",x"C4",x"00",x"BD",x"FB",
    x"F8",x"8E",x"C4",x"25",x"96",x"79",x"85",x"04",x"27",x"03",x"8E",x"C4",x"18",x"BD",x"FB",x"FE",
    x"8E",x"C3",x"E4",x"0D",x"79",x"2B",x"03",x"8E",x"C3",x"D0",x"C6",x"03",x"BD",x"FB",x"F8",x"C6",
    x"04",x"8E",x"C4",x"32",x"BD",x"FB",x"F8",x"86",x"24",x"7E",x"C1",x"2E",x"1B",x"7C",x"14",x"0C",
    x"1B",x"20",x"40",x"1B",x"20",x"58",x"1B",x"68",x"1F",x"10",x"16",x"1B",x"20",x"54",x"1F",x"12",
    x"14",x"1B",x"47",x"0D",x"0A",x"20",x"20",x"80",x"81",x"82",x"20",x"20",x"83",x"84",x"85",x"86",
    x"20",x"97",x"98",x"7E",x"7E",x"7E",x"99",x"9A",x"20",x"AB",x"7E",x"AC",x"AD",x"AE",x"AF",x"B0",
    x"0D",x"0A",x"20",x"20",x"87",x"88",x"20",x"89",x"20",x"8A",x"83",x"8B",x"8C",x"20",x"9B",x"9C",
    x"9D",x"7E",x"9E",x"9F",x"A0",x"20",x"87",x"B1",x"B2",x"5F",x"B3",x"B4",x"B5",x"0D",x"0A",x"20",
    x"20",x"87",x"7C",x"89",x"8D",x"83",x"8E",x"8A",x"8F",x"8C",x"20",x"87",x"7C",x"20",x"20",x"20",
    x"8F",x"8C",x"20",x"87",x"B6",x"B7",x"B8",x"B9",x"BA",x"BB",x"0D",x"0A",x"20",x"20",x"87",x"7C",
    x"8D",x"20",x"90",x"83",x"8E",x"8F",x"8C",x"20",x"A1",x"A2",x"A3",x"5F",x"A4",x"A5",x"A6",x"20",
    x"87",x"BC",x"20",x"20",x"BD",x"BE",x"8C",x"0D",x"0A",x"20",x"20",x"91",x"92",x"20",x"93",x"5F",
    x"94",x"20",x"95",x"96",x"20",x"A7",x"A8",x"5F",x"5F",x"5F",x"A9",x"AA",x"20",x"BF",x"C0",x"AD",
    x"AD",x"C1",x"C2",x"C3",x"20",x"1B",x"40",x"C4",x"C5",x"C6",x"C7",x"C8",x"C9",x"CA",x"CB",x"CC",
    x"CD",x"CE",x"1F",x"4E",x"5F",x"1B",x"44",x"1B",x"58",x"52",x"41",x"4D",x"3A",x"20",x"31",x"32",
    x"38",x"4B",x"0D",x"0A",x"04",x"42",x"41",x"53",x"49",x"43",x"20",x"31",x"32",x"38",x"20",x"4D",
    x"49",x"43",x"52",x"4F",x"53",x"4F",x"46",x"54",x"20",x"31",x"2E",x"30",x"0D",x"0A",x"04",x"42",
    x"41",x"53",x"49",x"43",x"20",x"4D",x"49",x"43",x"52",x"4F",x"53",x"4F",x"46",x"54",x"20",x"31",
    x"2E",x"30",x"0D",x"0A",x"04",x"52",x"16",x"42",x"65",x"73",x"65",x"61",x"75",x"0D",x"0A",x"04",
    x"52",x"16",x"42",x"65",x"67",x"6C",x"61",x"67",x"65",x"20",x"65",x"74",x"20",x"70",x"72",x"16",
    x"42",x"65",x"66",x"16",x"42",x"65",x"72",x"65",x"6E",x"63",x"65",x"73",x"0D",x"0A",x"04",x"1B",
    x"44",x"83",x"83",x"83",x"83",x"04",x"1B",x"58",x"0C",x"1F",x"44",x"41",x"1B",x"44",x"1B",x"57",
    x"20",x"20",x"66",x"65",x"6E",x"16",x"43",x"65",x"74",x"72",x"65",x"20",x"64",x"65",x"20",x"72",
    x"16",x"42",x"65",x"67",x"6C",x"61",x"67",x"65",x"20",x"64",x"75",x"20",x"63",x"72",x"61",x"79",
    x"6F",x"6E",x"20",x"6F",x"70",x"74",x"69",x"71",x"75",x"65",x"20",x"20",x"1B",x"56",x"18",x"0A",
    x"18",x"0A",x"18",x"0A",x"18",x"0A",x"18",x"0A",x"18",x"0A",x"1B",x"58",x"1F",x"4F",x"41",x"04",
    x"43",x"68",x"6F",x"69",x"73",x"69",x"72",x"20",x"73",x"61",x"20",x"70",x"61",x"6C",x"65",x"74",
    x"74",x"65",x"20",x"64",x"65",x"20",x"63",x"6F",x"75",x"6C",x"65",x"75",x"72",x"0D",x"0A",x"04",
    x"43",x"68",x"6F",x"69",x"73",x"69",x"72",x"20",x"6C",x"61",x"20",x"73",x"6F",x"75",x"72",x"69",
    x"73",x"0D",x"0A",x"04",x"43",x"68",x"6F",x"69",x"73",x"69",x"72",x"20",x"6C",x"65",x"20",x"63",
    x"72",x"61",x"79",x"6F",x"6E",x"20",x"6F",x"70",x"74",x"69",x"71",x"75",x"65",x"0D",x"0A",x"04",
    x"4D",x"65",x"74",x"74",x"72",x"65",x"20",x"6C",x"61",x"20",x"63",x"61",x"73",x"73",x"65",x"74",
    x"74",x"65",x"20",x"16",x"41",x"61",x"20",x"04",x"32",x"34",x"30",x"30",x"20",x"62",x"61",x"75",
    x"64",x"73",x"0D",x"0A",x"04",x"31",x"32",x"30",x"30",x"20",x"62",x"61",x"75",x"64",x"73",x"0D",
    x"0A",x"04",x"52",x"65",x"74",x"6F",x"75",x"72",x"20",x"16",x"41",x"61",x"20",x"6C",x"61",x"20",
    x"70",x"61",x"67",x"65",x"20",x"65",x"6E",x"2D",x"74",x"16",x"43",x"65",x"74",x"65",x"20",x"64",
    x"75",x"20",x"4D",x"4F",x"36",x"0D",x"0A",x"1B",x"44",x"83",x"83",x"83",x"83",x"04",x"80",x"80",
    x"80",x"80",x"80",x"80",x"80",x"FF",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"01",x"01",
    x"02",x"02",x"04",x"04",x"08",x"F0",x"02",x"02",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"80",x"80",x"40",x"3F",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"04",x"04",
    x"04",x"04",x"04",x"04",x"04",x"FC",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"11",x"11",
    x"12",x"12",x"14",x"14",x"18",x"18",x"10",x"10",x"20",x"20",x"40",x"40",x"80",x"80",x"20",x"20",
    x"10",x"10",x"08",x"08",x"04",x"04",x"20",x"20",x"20",x"20",x"A0",x"A0",x"60",x"60",x"04",x"04",
    x"04",x"04",x"04",x"04",x"04",x"04",x"01",x"01",x"02",x"02",x"04",x"04",x"08",x"08",x"00",x"00",
    x"00",x"00",x"80",x"80",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",
    x"00",x"30",x"48",x"48",x"84",x"84",x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"F0",x"10",
    x"10",x"10",x"10",x"10",x"10",x"10",x"1F",x"10",x"20",x"20",x"40",x"40",x"80",x"80",x"E0",x"20",
    x"10",x"10",x"08",x"08",x"04",x"04",x"3F",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"FC",x"04",
    x"04",x"04",x"04",x"04",x"04",x"04",x"20",x"20",x"10",x"08",x"04",x"03",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"C0",x"3F",x"00",x"00",x"00",x"00",x"00",x"03",x"0C",x"F0",x"10",x"10",
    x"20",x"40",x"80",x"00",x"00",x"00",x"80",x"80",x"80",x"80",x"80",x"80",x"40",x"40",x"10",x"10",
    x"08",x"08",x"04",x"02",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"7F",x"00",x"00",
    x"00",x"00",x"00",x"01",x"06",x"F8",x"20",x"20",x"40",x"40",x"80",x"00",x"00",x"00",x"04",x"04",
    x"04",x"04",x"04",x"04",x"08",x"08",x"40",x"40",x"80",x"80",x"80",x"80",x"80",x"80",x"00",x"01",
    x"02",x"04",x"08",x"08",x"10",x"10",x"7F",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"06",
    x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"40",x"20",x"20",x"08",x"08",
    x"04",x"04",x"04",x"04",x"04",x"04",x"00",x"00",x"03",x"04",x"08",x"10",x"20",x"20",x"3F",x"C0",
    x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"0C",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"80",x"40",x"20",x"10",x"10",x"40",x"40",x"20",x"10",x"08",x"04",x"03",x"00",x"7F",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"F8",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"FE",x"08",x"08",
    x"10",x"20",x"40",x"80",x"00",x"00",x"08",x"08",x"08",x"08",x"08",x"04",x"02",x"01",x"7F",x"00",
    x"00",x"00",x"00",x"00",x"00",x"80",x"FF",x"00",x"00",x"00",x"00",x"00",x"01",x"06",x"FC",x"00",
    x"00",x"00",x"7F",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"FC",x"04",x"04",x"04",x"02",x"01",
    x"00",x"08",x"0C",x"0C",x"0A",x"09",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"80",x"00",x"FF",
    x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"03",x"04",x"08",x"08",x"10",x"20",x"40",x"80",x"00",x"02",x"04",
    x"08",x"08",x"08",x"08",x"08",x"04",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",
    x"40",x"40",x"40",x"40",x"40",x"80",x"00",x"03",x"04",x"08",x"10",x"20",x"40",x"40",x"FF",x"00",
    x"00",x"00",x"00",x"00",x"00",x"01",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"FC",x"03",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"20",x"10",x"08",x"08",x"0E",x"0E",
    x"0E",x"0E",x"0E",x"0E",x"FF",x"FF",x"1C",x"1C",x"1C",x"1F",x"1F",x"1C",x"FC",x"FC",x"0E",x"0E",
    x"0E",x"FE",x"FE",x"0E",x"0E",x"0E",x"7F",x"FF",x"E0",x"E0",x"E0",x"E0",x"FF",x"7F",x"CE",x"EE",
    x"EE",x"EE",x"EF",x"EF",x"EF",x"CF",x"73",x"73",x"FB",x"FB",x"DF",x"8F",x"8F",x"07",x"9F",x"BF",
    x"80",x"9F",x"BF",x"B8",x"BF",x"9F",x"F1",x"FB",x"3B",x"FB",x"F3",x"03",x"FB",x"F1",x"FF",x"FF",
    x"83",x"83",x"83",x"83",x"FF",x"FF",x"38",x"B8",x"B8",x"B9",x"BB",x"BF",x"BE",x"3C",x"3C",x"7C",
    x"FC",x"DC",x"9C",x"1C",x"1C",x"1C",x"17",x"17",x"17",x"17",x"17",x"1F",x"00",x"00",x"01",x"0D",
    x"0D",x"0D",x"01",x"FF",x"00",x"00",x"08",x"08",x"08",x"08",x"08",x"F8",x"00",x"00",x"14",x"14",
    x"14",x"13",x"10",x"10",x"10",x"13",x"7E",x"00",x"00",x"FF",x"00",x"00",x"00",x"FE",x"48",x"48",
    x"48",x"88",x"08",x"08",x"08",x"08",x"00",x"00",x"1F",x"14",x"14",x"14",x"14",x"14",x"00",x"00",
    x"FF",x"00",x"FC",x"02",x"7C",x"80",x"00",x"00",x"F8",x"48",x"48",x"48",x"48",x"48",x"80",x"00",
    x"00",x"FF",x"00",x"00",x"00",x"FE",x"00",x"00",x"FF",x"00",x"FE",x"80",x"80",x"80",x"20",x"20",
    x"20",x"A8",x"70",x"20",x"00",x"00",x"04",x"04",x"04",x"15",x"0E",x"04",x"00",x"00",x"00",x"08",
    x"04",x"FE",x"FE",x"04",x"08",x"00",x"8C",x"8C",x"8F",x"8F",x"80",x"80",x"80",x"FF",x"00",x"00",
    x"FF",x"FF",x"00",x"00",x"00",x"FF",x"31",x"31",x"F1",x"F1",x"01",x"01",x"01",x"FF",x"8F",x"8C",
    x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"F1",x"31",x"31",x"31",x"31",x"31",x"31",x"31",x"FF",x"80",
    x"BF",x"A0",x"AA",x"95",x"88",x"87",x"FF",x"00",x"FF",x"00",x"AA",x"55",x"00",x"FF",x"FF",x"01",
    x"FD",x"05",x"A5",x"49",x"11",x"E1",x"8E",x"CE",x"95",x"BD",x"FB",x"FE",x"5F",x"34",x"04",x"4F",
    x"BD",x"CD",x"CC",x"30",x"02",x"8D",x"1F",x"BD",x"FB",x"FE",x"8D",x"1A",x"8D",x"28",x"A6",x"E4",
    x"8E",x"22",x"DA",x"48",x"EC",x"86",x"8D",x"16",x"8E",x"CE",x"84",x"BD",x"FB",x"FE",x"35",x"04",
    x"5C",x"C1",x"10",x"26",x"D8",x"39",x"C6",x"1B",x"3F",x"02",x"C6",x"7B",x"3F",x"82",x"84",x"0F",
    x"BD",x"CD",x"CC",x"7E",x"FB",x"FE",x"C6",x"20",x"3F",x"82",x"3F",x"04",x"8E",x"00",x"00",x"CE",
    x"CE",x"99",x"C6",x"05",x"A6",x"C0",x"A7",x"80",x"5A",x"26",x"FB",x"11",x"83",x"CE",x"A1",x"26",
    x"F1",x"8C",x"03",x"1F",x"23",x"E9",x"17",x"04",x"97",x"8E",x"00",x"00",x"CE",x"CE",x"A1",x"A6",
    x"C0",x"A7",x"80",x"11",x"83",x"CE",x"A6",x"26",x"F6",x"8C",x"03",x"1F",x"23",x"EE",x"39",x"8D",
    x"C9",x"8D",x"83",x"86",x"0E",x"B7",x"20",x"29",x"10",x"8E",x"00",x"2F",x"8E",x"00",x"43",x"31",
    x"A8",x"D1",x"1F",x"20",x"57",x"34",x"04",x"1F",x"10",x"E0",x"E0",x"1F",x"01",x"BF",x"20",x"32",
    x"34",x"10",x"1F",x"20",x"30",x"85",x"31",x"A8",x"30",x"10",x"BF",x"20",x"34",x"3F",x"0E",x"35",
    x"10",x"31",x"21",x"10",x"BF",x"20",x"34",x"3F",x"0E",x"10",x"8C",x"00",x"9F",x"23",x"CD",x"17",
    x"04",x"3E",x"CC",x"FF",x"FF",x"8E",x"07",x"94",x"ED",x"84",x"30",x"88",x"28",x"8C",x"19",x"3C",
    x"26",x"F6",x"86",x"7F",x"B7",x"00",x"15",x"CC",x"00",x"01",x"DD",x"BE",x"DD",x"C0",x"16",x"03",
    x"E7",x"BD",x"CC",x"BF",x"CE",x"21",x"00",x"8E",x"1A",x"40",x"10",x"8E",x"05",x"2E",x"17",x"04",
    x"0F",x"A6",x"84",x"6F",x"80",x"A7",x"C0",x"31",x"3F",x"26",x"F6",x"39",x"8E",x"21",x"00",x"CE",
    x"1A",x"40",x"8D",x"E6",x"CE",x"22",x"FA",x"86",x"0F",x"10",x"8E",x"00",x"00",x"8E",x"FF",x"FF",
    x"3F",x"3C",x"36",x"10",x"4A",x"2A",x"F6",x"39",x"86",x"22",x"1F",x"8B",x"BD",x"C1",x"20",x"8E",
    x"C6",x"D6",x"BF",x"20",x"70",x"8E",x"CD",x"FA",x"BD",x"FB",x"FE",x"7D",x"20",x"80",x"27",x"03",
    x"BD",x"FB",x"FE",x"8D",x"C7",x"10",x"CE",x"26",x"2C",x"03",x"B3",x"17",x"FF",x"41",x"4F",x"5F",
    x"BD",x"CA",x"53",x"B6",x"A7",x"E7",x"2A",x"FB",x"C6",x"0C",x"BD",x"FC",x"C7",x"86",x"0B",x"4A",
    x"26",x"FD",x"12",x"5A",x"26",x"F7",x"AC",x"01",x"8E",x"00",x"8C",x"30",x"1F",x"26",x"FC",x"8E",
    x"00",x"1E",x"CC",x"1E",x"A7",x"1F",x"9B",x"CE",x"A7",x"DC",x"36",x"10",x"97",x"DA",x"3D",x"3D",
    x"3D",x"3D",x"8E",x"E8",x"1C",x"CC",x"1B",x"2F",x"CE",x"A7",x"DC",x"36",x"10",x"97",x"DA",x"D7",
    x"DD",x"C6",x"22",x"1F",x"9B",x"1C",x"AF",x"D6",x"B3",x"2A",x"04",x"0C",x"B3",x"26",x"0F",x"58",
    x"CE",x"C9",x"DA",x"9E",x"BE",x"10",x"9E",x"C0",x"86",x"FF",x"97",x"B3",x"AD",x"D5",x"B6",x"A7",
    x"E7",x"2B",x"FB",x"1A",x"50",x"F6",x"A7",x"C3",x"2A",x"FB",x"F6",x"A7",x"C1",x"17",x"03",x"0F",
    x"8E",x"00",x"E8",x"30",x"1F",x"26",x"FC",x"96",x"D8",x"8A",x"20",x"B7",x"A7",x"DD",x"96",x"D8",
    x"48",x"AE",x"9F",x"22",x"D5",x"8D",x"0F",x"86",x"1C",x"9E",x"F6",x"8D",x"09",x"86",x"1E",x"9E",
    x"F8",x"8D",x"03",x"7E",x"C8",x"C3",x"B7",x"A7",x"DB",x"1F",x"10",x"F7",x"A7",x"DA",x"B7",x"A7",
    x"DA",x"39",x"10",x"CE",x"20",x"CC",x"BD",x"C8",x"61",x"3F",x"80",x"CC",x"00",x"FF",x"20",x"0D",
    x"CC",x"00",x"01",x"20",x"08",x"CC",x"01",x"00",x"20",x"03",x"CC",x"FF",x"00",x"9E",x"B6",x"30",
    x"86",x"10",x"9E",x"B8",x"31",x"A5",x"16",x"01",x"FD",x"17",x"03",x"D2",x"25",x"28",x"30",x"84",
    x"26",x"02",x"30",x"01",x"8C",x"01",x"3F",x"25",x"02",x"30",x"1F",x"9F",x"BE",x"10",x"8C",x"00",
    x"A7",x"25",x"04",x"10",x"8E",x"00",x"A6",x"10",x"9F",x"C0",x"17",x"04",x"10",x"24",x"07",x"8D",
    x"4B",x"24",x"03",x"D7",x"B3",x"39",x"86",x"0A",x"CE",x"C9",x"D8",x"E6",x"C2",x"F7",x"A7",x"C1",
    x"F6",x"A7",x"C1",x"2A",x"04",x"4A",x"26",x"F3",x"39",x"8B",x"05",x"97",x"B3",x"39",x"4C",x"5C",
    x"62",x"42",x"32",x"52",x"68",x"24",x"46",x"6E",x"C9",x"89",x"CB",x"86",x"CB",x"54",x"CA",x"45",
    x"C9",x"62",x"CC",x"C6",x"CC",x"AC",x"CB",x"41",x"CB",x"47",x"C9",x"6B",x"C9",x"70",x"C9",x"75",
    x"C9",x"7A",x"CA",x"3A",x"CC",x"AC",x"CC",x"C6",x"C9",x"62",x"C9",x"61",x"CE",x"CE",x"54",x"C6",
    x"05",x"10",x"AC",x"C4",x"23",x"0D",x"10",x"AC",x"42",x"22",x"08",x"AC",x"44",x"23",x"04",x"AC",
    x"46",x"23",x"07",x"33",x"48",x"5A",x"2A",x"E9",x"5F",x"39",x"1A",x"01",x"39",x"C6",x"18",x"8B",
    x"05",x"20",x"07",x"C6",x"05",x"3D",x"54",x"C3",x"04",x"02",x"34",x"06",x"C6",x"1F",x"3F",x"02",
    x"35",x"04",x"8D",x"02",x"35",x"04",x"CB",x"40",x"3F",x"82",x"C6",x"FC",x"D7",x"B3",x"D6",x"D8",
    x"5C",x"C4",x"0F",x"20",x"0C",x"31",x"A8",x"D8",x"1F",x"20",x"54",x"54",x"54",x"D1",x"D8",x"27",
    x"C9",x"96",x"D8",x"34",x"02",x"D7",x"D8",x"96",x"D8",x"48",x"8E",x"22",x"DA",x"30",x"86",x"9F",
    x"D5",x"A6",x"E4",x"8D",x"BE",x"17",x"FD",x"5E",x"96",x"D8",x"8D",x"B7",x"C6",x"8B",x"96",x"D8",
    x"44",x"C9",x"00",x"BD",x"FC",x"05",x"A6",x"E0",x"8D",x"A3",x"17",x"FD",x"49",x"96",x"D8",x"8D",
    x"9C",x"C6",x"8D",x"BD",x"FC",x"05",x"8E",x"CE",x"8D",x"BD",x"FB",x"FE",x"3F",x"04",x"D6",x"D8",
    x"1F",x"98",x"8E",x"03",x"20",x"ED",x"81",x"8C",x"04",x"FF",x"23",x"F9",x"EC",x"9F",x"22",x"D5",
    x"84",x"0F",x"97",x"D3",x"1F",x"98",x"C4",x"0F",x"D7",x"CF",x"44",x"44",x"44",x"44",x"97",x"D1",
    x"91",x"CF",x"24",x"02",x"96",x"CF",x"91",x"D3",x"24",x"02",x"96",x"D3",x"4C",x"34",x"02",x"8E",
    x"00",x"A8",x"10",x"9E",x"B4",x"BD",x"CC",x"8C",x"8D",x"6B",x"BD",x"CC",x"8C",x"10",x"9F",x"B4",
    x"96",x"CF",x"9B",x"D1",x"9B",x"D3",x"97",x"D4",x"26",x"0C",x"86",x"0F",x"97",x"CF",x"97",x"D1",
    x"97",x"D3",x"86",x"2D",x"97",x"D4",x"86",x"6C",x"97",x"CD",x"BD",x"CB",x"FD",x"86",x"03",x"97",
    x"D7",x"8E",x"22",x"CE",x"10",x"8E",x"22",x"C7",x"EC",x"81",x"ED",x"A1",x"0A",x"D7",x"26",x"F8",
    x"D6",x"C8",x"50",x"CB",x"6E",x"4F",x"1F",x"02",x"31",x"A8",x"30",x"D6",x"C8",x"54",x"DB",x"CC",
    x"CB",x"0E",x"1F",x"01",x"0D",x"D9",x"27",x"0E",x"34",x"30",x"9E",x"B6",x"10",x"9E",x"B8",x"BD",
    x"CC",x"8C",x"35",x"30",x"20",x"02",x"03",x"D9",x"BD",x"CC",x"8C",x"9F",x"B6",x"10",x"9F",x"B8",
    x"35",x"02",x"97",x"CD",x"39",x"C6",x"07",x"3D",x"C0",x"A4",x"50",x"1F",x"02",x"8E",x"00",x"A8",
    x"39",x"96",x"CD",x"4A",x"26",x"08",x"39",x"96",x"CD",x"4C",x"81",x"10",x"22",x"F8",x"C6",x"FC",
    x"D7",x"B3",x"8D",x"E1",x"34",x"20",x"31",x"A8",x"D0",x"86",x"07",x"97",x"B2",x"1F",x"20",x"BD",
    x"CC",x"25",x"53",x"C4",x"0F",x"5C",x"D7",x"B2",x"D7",x"CD",x"DC",x"C7",x"DD",x"CE",x"DC",x"C9",
    x"DD",x"D0",x"DC",x"CB",x"DD",x"D2",x"8E",x"00",x"A8",x"10",x"9E",x"B4",x"17",x"01",x"0D",x"35",
    x"20",x"10",x"9F",x"B4",x"20",x"45",x"10",x"8C",x"00",x"A0",x"24",x"05",x"3F",x"14",x"5D",x"2A",
    x"01",x"39",x"34",x"30",x"31",x"A8",x"D0",x"1F",x"20",x"C0",x"70",x"50",x"34",x"04",x"34",x"04",
    x"DD",x"C7",x"DD",x"CE",x"1F",x"10",x"C0",x"0B",x"67",x"E4",x"E0",x"E0",x"34",x"04",x"DD",x"D2",
    x"DD",x"CB",x"C6",x"70",x"E0",x"E0",x"E0",x"E0",x"DD",x"D0",x"DD",x"C9",x"9E",x"B6",x"10",x"9E",
    x"B8",x"17",x"00",x"C8",x"35",x"30",x"9F",x"B6",x"10",x"9F",x"B8",x"17",x"00",x"BE",x"8E",x"CE",
    x"88",x"BD",x"FB",x"FE",x"8D",x"17",x"D6",x"D1",x"58",x"58",x"58",x"58",x"DA",x"CF",x"A6",x"9F",
    x"22",x"D5",x"84",x"F0",x"9A",x"D3",x"ED",x"9F",x"22",x"D5",x"16",x"FB",x"D1",x"D6",x"C8",x"D1",
    x"CC",x"24",x"02",x"D6",x"CC",x"D1",x"CA",x"24",x"02",x"D6",x"CA",x"D7",x"D4",x"8E",x"22",x"CE",
    x"C6",x"03",x"D7",x"D7",x"EC",x"84",x"96",x"CD",x"3D",x"ED",x"81",x"0A",x"D7",x"26",x"F5",x"8E",
    x"22",x"CE",x"C6",x"03",x"D7",x"D7",x"96",x"D4",x"97",x"B2",x"EC",x"84",x"8D",x"07",x"ED",x"81",
    x"0A",x"D7",x"26",x"F2",x"39",x"6F",x"E2",x"34",x"06",x"4F",x"D6",x"B2",x"34",x"06",x"5F",x"E3",
    x"E4",x"6C",x"64",x"10",x"A3",x"62",x"25",x"F7",x"E6",x"64",x"4F",x"5A",x"32",x"65",x"39",x"8D",
    x"3F",x"9E",x"BA",x"10",x"9E",x"BC",x"8D",x"0A",x"9E",x"BE",x"10",x"9E",x"C0",x"9F",x"BA",x"10",
    x"9F",x"BC",x"30",x"1F",x"8D",x"0C",x"30",x"02",x"8D",x"08",x"30",x"1F",x"31",x"3F",x"8D",x"02",
    x"31",x"22",x"34",x"76",x"1F",x"20",x"86",x"28",x"3D",x"1E",x"01",x"44",x"56",x"54",x"54",x"30",
    x"8B",x"E6",x"63",x"C4",x"07",x"CE",x"F6",x"61",x"A6",x"C5",x"A8",x"84",x"A7",x"84",x"35",x"F6",
    x"34",x"02",x"B6",x"A7",x"C0",x"8A",x"01",x"B7",x"A7",x"C0",x"35",x"82",x"8D",x"F2",x"20",x"D2",
    x"B7",x"A7",x"C0",x"A6",x"62",x"10",x"3F",x"B6",x"A7",x"C0",x"8A",x"20",x"B7",x"A7",x"C0",x"39",
    x"50",x"41",x"4C",x"45",x"54",x"54",x"45",x"20",x"43",x"46",x"47",x"00",x"7D",x"20",x"80",x"27",
    x"EE",x"1F",x"43",x"4F",x"8D",x"19",x"8D",x"07",x"BD",x"C7",x"86",x"5F",x"7E",x"CA",x"51",x"86",
    x"FF",x"8E",x"22",x"DA",x"3F",x"BC",x"7D",x"20",x"80",x"27",x"D4",x"1F",x"43",x"86",x"FF",x"34",
    x"02",x"7F",x"20",x"49",x"C6",x"10",x"10",x"8E",x"22",x"FA",x"8E",x"CC",x"90",x"8D",x"58",x"5F",
    x"8D",x"47",x"8E",x"23",x"0A",x"BF",x"21",x"97",x"8E",x"24",x"0A",x"BF",x"21",x"99",x"8E",x"24",
    x"B0",x"86",x"01",x"10",x"8E",x"00",x"01",x"C6",x"02",x"8D",x"2E",x"C6",x"0C",x"8E",x"CC",x"A0",
    x"10",x"8E",x"22",x"4F",x"8D",x"31",x"8E",x"02",x"00",x"9F",x"4C",x"CC",x"00",x"20",x"DD",x"47",
    x"CC",x"22",x"DA",x"DD",x"AA",x"CC",x"40",x"03",x"97",x"4B",x"8D",x"0D",x"35",x"02",x"97",x"49",
    x"8E",x"00",x"01",x"C6",x"07",x"8D",x"02",x"C6",x"06",x"34",x"02",x"B6",x"A7",x"C0",x"84",x"DF",
    x"9D",x"FA",x"5D",x"26",x"0A",x"35",x"82",x"A6",x"80",x"A7",x"A0",x"5A",x"26",x"F9",x"39",x"86",
    x"20",x"B7",x"A7",x"DD",x"8E",x"00",x"00",x"BD",x"F4",x"75",x"86",x"2F",x"B7",x"A7",x"DD",x"BD",
    x"F4",x"75",x"3F",x"0A",x"5D",x"26",x"04",x"3F",x"16",x"24",x"E4",x"1F",x"34",x"39",x"7D",x"20",
    x"79",x"2A",x"2A",x"34",x"06",x"BE",x"20",x"7A",x"10",x"BE",x"20",x"7C",x"F6",x"20",x"E3",x"BD",
    x"F0",x"AE",x"30",x"8B",x"F6",x"20",x"E4",x"BD",x"F0",x"AE",x"31",x"AB",x"BF",x"20",x"7A",x"10",
    x"BF",x"20",x"7C",x"7F",x"20",x"E3",x"7F",x"20",x"E4",x"3F",x"40",x"35",x"86",x"34",x"7F",x"86",
    x"20",x"1F",x"8B",x"8D",x"04",x"32",x"61",x"35",x"FE",x"1A",x"50",x"BE",x"20",x"67",x"34",x"18",
    x"CE",x"A7",x"C0",x"8E",x"F9",x"3B",x"BF",x"20",x"67",x"86",x"A7",x"1F",x"8B",x"10",x"8E",x"20",
    x"CD",x"86",x"FF",x"A7",x"42",x"6D",x"C4",x"8E",x"04",x"00",x"7E",x"F8",x"54",x"7D",x"20",x"79",
    x"2A",x"02",x"3F",x"BE",x"B6",x"A7",x"C0",x"84",x"02",x"8B",x"FF",x"39",x"8E",x"22",x"C2",x"34",
    x"56",x"CE",x"CD",x"F2",x"86",x"2F",x"A7",x"84",x"EC",x"E4",x"6C",x"84",x"ED",x"E4",x"A3",x"C4",
    x"24",x"F8",x"33",x"42",x"30",x"01",x"11",x"83",x"CD",x"FA",x"26",x"E8",x"86",x"04",x"A7",x"84",
    x"35",x"D6",x"03",x"E8",x"00",x"64",x"00",x"0A",x"00",x"01",x"1B",x"4E",x"1B",x"5F",x"0C",x"1F",
    x"22",x"21",x"1B",x"4F",x"0C",x"1B",x"4E",x"1F",x"20",x"20",x"1F",x"45",x"49",x"52",x"1F",x"53",
    x"41",x"56",x"1F",x"53",x"51",x"42",x"1F",x"52",x"62",x"8E",x"8F",x"90",x"0A",x"08",x"08",x"08",
    x"91",x"5F",x"92",x"0A",x"08",x"08",x"08",x"93",x"94",x"95",x"04",x"1F",x"46",x"62",x"80",x"81",
    x"82",x"0A",x"08",x"08",x"08",x"83",x"89",x"85",x"0A",x"08",x"08",x"08",x"86",x"8A",x"88",x"1F",
    x"4C",x"62",x"80",x"81",x"82",x"0A",x"08",x"08",x"08",x"83",x"84",x"85",x"0A",x"08",x"08",x"08",
    x"86",x"87",x"88",x"04",x"00",x"30",x"00",x"48",x"01",x"08",x"01",x"20",x"00",x"60",x"00",x"78",
    x"01",x"08",x"01",x"20",x"00",x"90",x"00",x"A8",x"01",x"08",x"01",x"20",x"00",x"28",x"00",x"A7",
    x"00",x"C0",x"00",x"CF",x"00",x"30",x"00",x"A0",x"00",x"A0",x"00",x"B0",x"00",x"30",x"00",x"A0",
    x"00",x"0B",x"00",x"7B",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"04",x"09",x"09",x"09",
    x"09",x"09",x"09",x"09",x"04",x"1F",x"45",x"59",x"04",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",
    x"EF",x"FF",x"FF",x"F0",x"00",x"00",x"34",x"46",x"CE",x"A7",x"CC",x"EC",x"42",x"84",x"3F",x"81",
    x"14",x"26",x"08",x"A6",x"42",x"85",x"C0",x"26",x"36",x"35",x"C6",x"C4",x"FB",x"86",x"14",x"ED",
    x"42",x"A6",x"41",x"8A",x"01",x"A7",x"41",x"CA",x"04",x"E7",x"43",x"A6",x"41",x"8A",x"01",x"A7",
    x"41",x"EC",x"C4",x"43",x"85",x"0C",x"26",x"17",x"53",x"C5",x"44",x"26",x"12",x"A6",x"43",x"84",
    x"FB",x"A7",x"43",x"E6",x"41",x"C4",x"FE",x"E7",x"41",x"8A",x"04",x"A7",x"43",x"35",x"C6",x"96",
    x"79",x"8A",x"C0",x"97",x"79",x"86",x"1F",x"A7",x"42",x"20",x"E2",x"0F",x"2B",x"C6",x"0C",x"3F",
    x"02",x"C6",x"1B",x"3F",x"02",x"C6",x"68",x"3F",x"02",x"8D",x"09",x"3F",x"0A",x"C1",x"20",x"26",
    x"FA",x"7E",x"C0",x"00",x"8E",x"D0",x"00",x"3F",x"06",x"8D",x"03",x"7A",x"A7",x"C0",x"CE",x"00",
    x"00",x"CC",x"28",x"C8",x"34",x"46",x"E6",x"80",x"27",x"08",x"A6",x"80",x"8D",x"12",x"26",x"FC",
    x"20",x"F4",x"E6",x"80",x"27",x"08",x"A6",x"80",x"8D",x"06",x"26",x"FA",x"20",x"E8",x"35",x"C6",
    x"A7",x"C4",x"33",x"C8",x"28",x"6A",x"63",x"26",x"10",x"34",x"02",x"6A",x"63",x"86",x"C8",x"A7",
    x"64",x"EE",x"65",x"33",x"41",x"EF",x"65",x"35",x"02",x"5A",x"39",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"08",x"00",x"00",x"01",x"FF",x"2A",x"80",x"03",x"81",x"00",x"03",x"83",x"85",x"81",x"02",x"95",
    x"00",x"04",x"AF",x"AB",x"BF",x"AF",x"03",x"FF",x"00",x"03",x"BF",x"FF",x"BF",x"29",x"FF",x"00",
    x"01",x"BF",x"02",x"FF",x"00",x"05",x"DF",x"D7",x"AF",x"8B",x"85",x"02",x"81",x"00",x"06",x"85",
    x"81",x"83",x"85",x"83",x"95",x"02",x"81",x"00",x"0F",x"A8",x"C2",x"A1",x"85",x"9D",x"DC",x"94",
    x"9E",x"8A",x"87",x"80",x"81",x"87",x"DF",x"BF",x"0D",x"FF",x"00",x"01",x"AA",x"05",x"FF",x"00",
    x"01",x"BF",x"0F",x"FF",x"00",x"01",x"AF",x"03",x"FF",x"00",x"0F",x"D5",x"FF",x"AA",x"FF",x"AF",
    x"BF",x"DD",x"DF",x"AA",x"AB",x"AA",x"BD",x"F7",x"FD",x"95",x"02",x"8A",x"0A",x"FF",x"29",x"00",
    x"00",x"09",x"03",x"57",x"3F",x"FF",x"D7",x"FF",x"57",x"DF",x"BF",x"03",x"FF",x"00",x"01",x"DF",
    x"37",x"FF",x"00",x"01",x"7F",x"06",x"FF",x"00",x"01",x"FE",x"02",x"7F",x"00",x"02",x"FF",x"7F",
    x"02",x"FF",x"00",x"05",x"7F",x"FF",x"3F",x"5F",x"17",x"11",x"FF",x"00",x"01",x"FE",x"03",x"FF",
    x"00",x"01",x"DF",x"05",x"FF",x"00",x"03",x"FD",x"FF",x"D5",x"03",x"FF",x"00",x"01",x"FD",x"03",
    x"FF",x"00",x"01",x"EF",x"03",x"FF",x"00",x"03",x"F7",x"FF",x"57",x"04",x"FF",x"00",x"09",x"7F",
    x"55",x"FF",x"AA",x"F7",x"FF",x"5F",x"5D",x"7F",x"02",x"D5",x"00",x"03",x"BD",x"55",x"5D",x"0A",
    x"FF",x"11",x"00",x"00",x"04",x"01",x"00",x"02",x"04",x"05",x"00",x"00",x"01",x"04",x"02",x"00",
    x"00",x"09",x"01",x"03",x"15",x"01",x"02",x"05",x"2F",x"0F",x"3F",x"02",x"7F",x"00",x"03",x"F7",
    x"FF",x"57",x"49",x"FF",x"00",x"03",x"7F",x"FF",x"7F",x"07",x"FF",x"00",x"01",x"7F",x"11",x"FF",
    x"00",x"01",x"57",x"07",x"FF",x"00",x"03",x"5F",x"FF",x"7F",x"03",x"FF",x"00",x"01",x"7F",x"15",
    x"FF",x"00",x"01",x"7F",x"13",x"FF",x"0E",x"00",x"00",x"02",x"0A",x"7B",x"02",x"80",x"04",x"00",
    x"00",x"01",x"02",x"02",x"00",x"00",x"09",x"07",x"0F",x"57",x"7B",x"FF",x"AF",x"FF",x"5F",x"7F",
    x"2C",x"FF",x"00",x"1A",x"FE",x"FF",x"FE",x"FF",x"FE",x"FF",x"F8",x"FA",x"F4",x"FD",x"FA",x"FC",
    x"EA",x"FA",x"E0",x"FD",x"F0",x"F4",x"F8",x"FA",x"F0",x"FA",x"FC",x"FF",x"FC",x"FF",x"02",x"FE",
    x"06",x"FF",x"00",x"02",x"FA",x"FB",x"12",x"FF",x"00",x"01",x"FE",x"05",x"FF",x"00",x"08",x"FE",
    x"FF",x"FA",x"FF",x"FE",x"FD",x"FA",x"FF",x"02",x"FA",x"00",x"2A",x"F4",x"FD",x"FA",x"F7",x"EA",
    x"FA",x"E8",x"FD",x"D0",x"F5",x"EA",x"FE",x"EA",x"FA",x"D5",x"F5",x"FA",x"FF",x"EA",x"FE",x"D5",
    x"FD",x"E8",x"FF",x"FB",x"FF",x"E8",x"FD",x"D5",x"F5",x"EA",x"FF",x"FA",x"FB",x"D5",x"F5",x"F7",
    x"F5",x"FA",x"FF",x"AA",x"FD",x"0A",x"FF",x"0E",x"00",x"00",x"0C",x"5E",x"3E",x"0A",x"00",x"AB",
    x"02",x"BF",x"5F",x"7F",x"AA",x"FF",x"AA",x"0D",x"FF",x"00",x"01",x"AB",x"05",x"FF",x"00",x"01",
    x"FE",x"13",x"FF",x"00",x"06",x"FA",x"FF",x"EF",x"FF",x"F5",x"FA",x"02",x"EA",x"00",x"0E",x"AA",
    x"BF",x"97",x"FF",x"AB",x"FF",x"AA",x"A9",x"A0",x"B5",x"05",x"2B",x"0A",x"AA",x"13",x"00",x"00",
    x"01",x"80",x"03",x"00",x"00",x"41",x"80",x"00",x"A0",x"80",x"A0",x"80",x"A0",x"80",x"D0",x"A0",
    x"E8",x"80",x"AD",x"80",x"D5",x"94",x"EA",x"80",x"AD",x"80",x"A5",x"20",x"51",x"A8",x"AA",x"8A",
    x"AD",x"15",x"95",x"02",x"AA",x"00",x"A9",x"80",x"B5",x"11",x"AA",x"A8",x"AA",x"02",x"A5",x"00",
    x"4A",x"00",x"A0",x"00",x"A1",x"00",x"81",x"00",x"AA",x"00",x"A8",x"08",x"85",x"00",x"48",x"80",
    x"AA",x"A0",x"A8",x"80",x"B5",x"00",x"E8",x"02",x"AA",x"00",x"05",x"A0",x"B5",x"00",x"5A",x"A8",
    x"04",x"AA",x"00",x"04",x"7E",x"AA",x"FA",x"AA",x"0A",x"FF",x"0C",x"00",x"00",x"01",x"02",x"02",
    x"00",x"00",x"0B",x"AA",x"F5",x"14",x"FF",x"78",x"FD",x"AA",x"F5",x"BE",x"FF",x"F7",x"14",x"FF",
    x"00",x"02",x"7F",x"BF",x"0D",x"FF",x"00",x"01",x"FE",x"04",x"FF",x"00",x"06",x"DF",x"55",x"FD",
    x"AE",x"F5",x"7D",x"02",x"7F",x"03",x"FF",x"00",x"05",x"FE",x"D5",x"55",x"5F",x"57",x"03",x"FF",
    x"00",x"07",x"FD",x"FF",x"55",x"0F",x"00",x"05",x"00",x"02",x"05",x"00",x"01",x"1A",x"17",x"00",
    x"00",x"2B",x"01",x"00",x"04",x"10",x"18",x"00",x"10",x"00",x"51",x"00",x"50",x"01",x"2A",x"00",
    x"50",x"00",x"50",x"55",x"4B",x"02",x"B5",x"A8",x"55",x"04",x"52",x"54",x"B5",x"20",x"F5",x"AE",
    x"5F",x"15",x"4F",x"02",x"15",x"00",x"55",x"00",x"43",x"00",x"05",x"00",x"05",x"03",x"00",x"00",
    x"1A",x"0A",x"80",x"50",x"00",x"15",x"00",x"42",x"00",x"14",x"00",x"01",x"00",x"40",x"10",x"80",
    x"00",x"01",x"00",x"55",x"00",x"42",x"82",x"B5",x"80",x"54",x"00",x"0A",x"FF",x"09",x"00",x"00",
    x"0E",x"03",x"02",x"5F",x"15",x"AB",x"55",x"BF",x"AA",x"5F",x"BF",x"7F",x"FD",x"FF",x"77",x"03",
    x"FF",x"00",x"01",x"F7",x"23",x"FF",x"00",x"03",x"7F",x"FF",x"7F",x"02",x"FF",x"00",x"04",x"FB",
    x"55",x"EA",x"57",x"05",x"FF",x"00",x"04",x"5F",x"AF",x"47",x"BD",x"03",x"FF",x"00",x"0E",x"FA",
    x"FC",x"FD",x"FB",x"FF",x"D5",x"EA",x"01",x"AA",x"57",x"7F",x"05",x"0A",x"04",x"12",x"00",x"00",
    x"03",x"20",x"00",x"80",x"05",x"00",x"00",x"43",x"20",x"00",x"A1",x"00",x"BC",x"3E",x"7F",x"55",
    x"AE",x"14",x"AA",x"0A",x"95",x"04",x"28",x"00",x"A8",x"51",x"AD",x"11",x"2A",x"10",x"AA",x"40",
    x"A5",x"80",x"5A",x"50",x"EA",x"50",x"AA",x"51",x"5F",x"55",x"6B",x"15",x"AA",x"15",x"56",x"00",
    x"02",x"04",x"AA",x"10",x"AA",x"11",x"57",x"05",x"2A",x"15",x"2A",x"13",x"AF",x"00",x"0A",x"05",
    x"AA",x"15",x"A8",x"11",x"5B",x"15",x"2A",x"55",x"AA",x"15",x"57",x"0A",x"FF",x"09",x"00",x"00",
    x"0C",x"A0",x"55",x"BD",x"55",x"FD",x"EA",x"DF",x"F5",x"FF",x"7F",x"FF",x"7F",x"03",x"FF",x"00",
    x"03",x"DF",x"FF",x"7F",x"25",x"FF",x"00",x"01",x"FA",x"05",x"FF",x"00",x"03",x"EA",x"AF",x"55",
    x"05",x"FF",x"00",x"03",x"5F",x"BF",x"57",x"04",x"FF",x"00",x"0B",x"BF",x"5F",x"FF",x"57",x"FD",
    x"FA",x"AF",x"55",x"BD",x"50",x"D5",x"0D",x"00",x"00",x"01",x"40",x"04",x"00",x"00",x"02",x"01",
    x"05",x"02",x"01",x"05",x"00",x"00",x"07",x"11",x"00",x"40",x"00",x"04",x"01",x"FD",x"02",x"FF",
    x"00",x"3A",x"AB",x"57",x"05",x"95",x"02",x"55",x"0B",x"57",x"55",x"BD",x"05",x"95",x"03",x"53",
    x"00",x"80",x"00",x"05",x"00",x"51",x"02",x"46",x"40",x"BD",x"55",x"FD",x"FB",x"F7",x"FB",x"BF",
    x"55",x"BD",x"1F",x"55",x"0B",x"57",x"15",x"BD",x"54",x"F5",x"EA",x"55",x"F5",x"AF",x"55",x"FD",
    x"55",x"F5",x"AA",x"AD",x"45",x"AD",x"55",x"F5",x"3A",x"57",x"D5",x"AF",x"0A",x"FF",x"09",x"00",
    x"00",x"06",x"0B",x"FF",x"FE",x"AF",x"57",x"5F",x"02",x"FF",x"00",x"01",x"FB",x"31",x"FF",x"00",
    x"14",x"AA",x"FF",x"EA",x"5A",x"A8",x"EA",x"A8",x"EA",x"D5",x"FF",x"FA",x"FF",x"FA",x"FF",x"AE",
    x"FF",x"F6",x"5E",x"A8",x"EA",x"02",x"A8",x"00",x"06",x"A0",x"78",x"00",x"40",x"00",x"80",x"11",
    x"00",x"00",x"0B",x"42",x"E2",x"FA",x"AA",x"AB",x"AF",x"5F",x"0A",x"2A",x"02",x"21",x"05",x"00",
    x"00",x"02",x"F8",x"AA",x"03",x"FF",x"00",x"0E",x"AF",x"6A",x"AA",x"FE",x"A4",x"AD",x"7F",x"FF",
    x"AA",x"FB",x"AA",x"AF",x"02",x"1E",x"03",x"00",x"00",x"01",x"80",x"03",x"00",x"02",x"AA",x"00",
    x"0B",x"FA",x"AA",x"57",x"5F",x"FF",x"FA",x"FF",x"AA",x"FD",x"57",x"5F",x"02",x"EA",x"00",x"0E",
    x"A8",x"AA",x"44",x"52",x"40",x"56",x"FA",x"EA",x"AA",x"AB",x"50",x"5E",x"00",x"4A",x"02",x"AA",
    x"00",x"05",x"A0",x"54",x"40",x"5E",x"AA",x"0A",x"FF",x"05",x"00",x"00",x"05",x"07",x"0F",x"2B",
    x"AF",x"AA",x"02",x"FF",x"00",x"04",x"AF",x"FB",x"BF",x"AE",x"03",x"FF",x"00",x"03",x"FB",x"FF",
    x"EA",x"13",x"FF",x"00",x"01",x"FE",x"19",x"FF",x"00",x"10",x"55",x"AF",x"AA",x"D5",x"04",x"15",
    x"54",x"57",x"AA",x"BF",x"AA",x"FF",x"F5",x"D7",x"AA",x"A1",x"1D",x"00",x"02",x"80",x"00",x"07",
    x"C1",x"E3",x"EF",x"AA",x"AD",x"A8",x"D7",x"02",x"50",x"00",x"02",x"00",x"20",x"05",x"00",x"00",
    x"02",x"E8",x"AA",x"02",x"FF",x"00",x"0D",x"F8",x"00",x"40",x"A8",x"A9",x"00",x"FD",x"FE",x"FF",
    x"EA",x"AB",x"A8",x"B4",x"09",x"00",x"02",x"A8",x"00",x"04",x"EA",x"AA",x"FD",x"FE",x"02",x"FF",
    x"00",x"16",x"EA",x"AA",x"B5",x"A0",x"D5",x"88",x"A8",x"02",x"A8",x"AA",x"B5",x"80",x"D5",x"03",
    x"A8",x"20",x"AD",x"00",x"B4",x"80",x"A8",x"00",x"02",x"A0",x"00",x"02",x"B5",x"80",x"0A",x"FF",
    x"02",x"00",x"00",x"11",x"0A",x"75",x"A0",x"DF",x"BD",x"7A",x"FF",x"FD",x"AA",x"FF",x"AA",x"FF",
    x"D7",x"EF",x"AA",x"FF",x"BF",x"09",x"FF",x"00",x"03",x"D5",x"FF",x"FA",x"03",x"FF",x"00",x"03",
    x"F7",x"FF",x"FD",x"05",x"FF",x"00",x"03",x"7F",x"FF",x"BF",x"03",x"FF",x"00",x"01",x"D7",x"0E",
    x"FF",x"00",x"1C",x"FE",x"F7",x"FF",x"F4",x"50",x"40",x"E8",x"00",x"50",x"00",x"57",x"55",x"5F",
    x"55",x"FF",x"AF",x"FF",x"AE",x"5F",x"15",x"2F",x"15",x"2B",x"01",x"03",x"00",x"03",x"05",x"17",
    x"00",x"00",x"04",x"E8",x"F0",x"E0",x"40",x"0B",x"00",x"00",x"04",x"7A",x"1D",x"7F",x"F5",x"04",
    x"00",x"00",x"08",x"40",x"00",x"20",x"40",x"50",x"80",x"50",x"80",x"0A",x"00",x"00",x"23",x"50",
    x"20",x"5A",x"84",x"6A",x"55",x"F5",x"A8",x"54",x"15",x"6A",x"00",x"D5",x"02",x"51",x"A0",x"52",
    x"04",x"22",x"A8",x"54",x"00",x"50",x"80",x"6A",x"01",x"0A",x"02",x"55",x"07",x"57",x"1F",x"7F",
    x"2A",x"7F",x"0A",x"FF",x"00",x"0F",x"00",x"0A",x"80",x"A8",x"55",x"AD",x"55",x"7F",x"BE",x"AA",
    x"55",x"AF",x"55",x"FF",x"BE",x"03",x"FF",x"00",x"01",x"F7",x"0D",x"FF",x"00",x"05",x"77",x"FF",
    x"7F",x"FF",x"FD",x"19",x"FF",x"00",x"08",x"FB",x"FF",x"55",x"AF",x"57",x"95",x"00",x"05",x"02",
    x"00",x"00",x"03",x"11",x"AF",x"7F",x"04",x"FF",x"00",x"04",x"EE",x"55",x"FF",x"7F",x"03",x"FF",
    x"00",x"09",x"D7",x"EF",x"55",x"F5",x"78",x"FA",x"00",x"2A",x"05",x"22",x"00",x"00",x"04",x"0D",
    x"7D",x"FD",x"80",x"16",x"00",x"00",x"18",x"02",x"00",x"15",x"50",x"D4",x"C4",x"A8",x"40",x"A5",
    x"00",x"81",x"00",x"A0",x"00",x"A0",x"45",x"05",x"07",x"57",x"07",x"AF",x"15",x"AF",x"57",x"02",
    x"BF",x"03",x"FF",x"00",x"06",x"5F",x"FE",x"7C",x"FE",x"FC",x"F8",x"0A",x"FF",x"00",x"0B",x"00",
    x"80",x"40",x"00",x"A5",x"05",x"F5",x"55",x"57",x"53",x"FF",x"02",x"FD",x"00",x"10",x"D5",x"F7",
    x"7F",x"FF",x"FB",x"FF",x"D5",x"F7",x"57",x"FF",x"FB",x"FF",x"EB",x"FF",x"5F",x"FD",x"02",x"FF",
    x"00",x"09",x"EA",x"FF",x"AA",x"FF",x"F7",x"FF",x"FB",x"FF",x"FB",x"15",x"FF",x"00",x"01",x"7F",
    x"03",x"FF",x"00",x"04",x"BF",x"FF",x"55",x"D5",x"03",x"00",x"00",x"02",x"5A",x"FA",x"03",x"FF",
    x"00",x"05",x"FB",x"52",x"00",x"EA",x"F5",x"02",x"FF",x"00",x"07",x"F3",x"F0",x"F8",x"E0",x"F0",
    x"00",x"D4",x"03",x"00",x"00",x"01",x"68",x"23",x"00",x"00",x"01",x"C0",x"11",x"00",x"02",x"03",
    x"00",x"03",x"0B",x"11",x"57",x"02",x"47",x"02",x"0F",x"00",x"0A",x"0E",x"1F",x"0F",x"5F",x"1F",
    x"7F",x"3E",x"3F",x"5D",x"7F",x"02",x"7C",x"00",x"02",x"FC",x"FF",x"06",x"FC",x"00",x"04",x"E8",
    x"E0",x"D0",x"F0",x"02",x"C0",x"07",x"00",x"0A",x"FF",x"07",x"00",x"00",x"11",x"40",x"A8",x"A0",
    x"7C",x"5F",x"FF",x"FE",x"BF",x"AA",x"FF",x"5F",x"FF",x"FB",x"FF",x"AE",x"EF",x"AF",x"03",x"FF",
    x"00",x"03",x"FB",x"FF",x"EA",x"05",x"FF",x"00",x"01",x"EA",x"0D",x"FF",x"00",x"01",x"FE",x"05",
    x"FF",x"00",x"01",x"AF",x"05",x"FF",x"00",x"01",x"FE",x"03",x"FF",x"00",x"04",x"FD",x"FC",x"F0",
    x"80",x"05",x"00",x"00",x"0F",x"E8",x"AA",x"FE",x"AE",x"FF",x"05",x"0A",x"00",x"E0",x"A0",x"F8",
    x"E8",x"FC",x"7E",x"2A",x"2F",x"00",x"00",x"01",x"02",x"03",x"03",x"03",x"0F",x"00",x"01",x"1F",
    x"02",x"3F",x"00",x"09",x"FF",x"FB",x"FF",x"57",x"FB",x"D3",x"EA",x"A2",x"A5",x"02",x"C0",x"00",
    x"02",x"40",x"00",x"02",x"80",x"1D",x"00",x"0A",x"FF",x"0C",x"00",x"00",x"0D",x"80",x"C0",x"F0",
    x"F8",x"AA",x"FD",x"AE",x"DF",x"57",x"5F",x"EA",x"FD",x"EA",x"02",x"FD",x"00",x"04",x"FF",x"F5",
    x"FF",x"BF",x"05",x"FF",x"00",x"03",x"D5",x"FF",x"EA",x"13",x"FF",x"00",x"01",x"BF",x"03",x"FF",
    x"00",x"05",x"F5",x"E5",x"EF",x"17",x"00",x"02",x"01",x"08",x"00",x"00",x"05",x"C0",x"E0",x"F0",
    x"A0",x"40",x"15",x"00",x"00",x"01",x"01",x"03",x"00",x"00",x"0A",x"01",x"00",x"01",x"02",x"03",
    x"00",x"05",x"02",x"05",x"08",x"02",x"1F",x"02",x"0F",x"00",x"05",x"1F",x"0F",x"1F",x"3F",x"5F",
    x"03",x"3F",x"03",x"7F",x"0A",x"FF",x"00",x"03",x"FE",x"FF",x"FE",x"05",x"FF",x"00",x"08",x"FE",
    x"FF",x"FD",x"AF",x"AA",x"BD",x"AA",x"55",x"20",x"00",x"0A",x"FF",x"14",x"00",x"00",x"13",x"80",
    x"00",x"80",x"C0",x"40",x"A0",x"00",x"BC",x"A0",x"FA",x"F5",x"EB",x"D5",x"FF",x"DF",x"FE",x"FD",
    x"FF",x"55",x"05",x"FF",x"00",x"03",x"F5",x"FF",x"D7",x"05",x"FF",x"00",x"01",x"FD",x"0F",x"FF",
    x"02",x"7F",x"00",x"01",x"FF",x"02",x"7F",x"00",x"04",x"BF",x"5F",x"BF",x"3F",x"02",x"7F",x"00",
    x"04",x"2F",x"5F",x"2F",x"3F",x"04",x"1F",x"00",x"04",x"2F",x"17",x"3F",x"0B",x"03",x"0F",x"00",
    x"07",x"1F",x"2F",x"17",x"1F",x"2F",x"5F",x"3F",x"02",x"7F",x"00",x"0A",x"FF",x"BF",x"7F",x"BF",
    x"7F",x"BF",x"EF",x"8B",x"5F",x"AB",x"02",x"5F",x"00",x"02",x"BF",x"7F",x"15",x"FF",x"00",x"02",
    x"EA",x"F2",x"02",x"E0",x"02",x"80",x"00",x"01",x"00",x"02",x"80",x"00",x"02",x"C0",x"80",x"02",
    x"C0",x"00",x"09",x"E0",x"A0",x"D8",x"A8",x"EA",x"45",x"A2",x"80",x"50",x"11",x"00",x"00",x"01",
    x"02",x"02",x"01",x"00",x"06",x"02",x"07",x"00",x"0A",x"04",x"28",x"03",x"00",x"00",x"01",x"10",
    x"0A",x"FF",x"1E",x"00",x"00",x"0A",x"A0",x"50",x"F8",x"5C",x"DE",x"BE",x"7F",x"55",x"FF",x"7F",
    x"03",x"FF",x"00",x"03",x"EB",x"FF",x"57",x"03",x"FF",x"00",x"03",x"BB",x"FF",x"77",x"35",x"FF",
    x"00",x"01",x"D7",x"11",x"FF",x"00",x"04",x"FD",x"FF",x"FC",x"FE",x"02",x"FC",x"02",x"F8",x"02",
    x"F0",x"02",x"E0",x"00",x"04",x"C0",x"04",x"00",x"40",x"0F",x"00",x"00",x"13",x"A0",x"F0",x"BD",
    x"55",x"F5",x"58",x"2A",x"54",x"2A",x"10",x"05",x"00",x"15",x"01",x"22",x"05",x"01",x"00",x"04",
    x"03",x"00",x"00",x"0B",x"A0",x"00",x"80",x"01",x"05",x"01",x"0A",x"04",x"08",x"00",x"20",x"03",
    x"40",x"0A",x"FF",x"26",x"00",x"02",x"80",x"02",x"C0",x"00",x"03",x"F0",x"C0",x"F0",x"03",x"E0",
    x"02",x"F0",x"00",x"04",x"F8",x"F0",x"F8",x"EA",x"07",x"FF",x"00",x"01",x"FE",x"2F",x"FF",x"02",
    x"FE",x"04",x"FF",x"02",x"F8",x"00",x"05",x"F0",x"FC",x"D4",x"D7",x"40",x"02",x"00",x"00",x"03",
    x"80",x"00",x"50",x"03",x"00",x"00",x"01",x"80",x"1A",x"00",x"00",x"03",x"C0",x"E8",x"40",x"03",
    x"50",x"00",x"06",x"00",x"60",x"40",x"E0",x"40",x"C0",x"04",x"00",x"00",x"08",x"01",x"05",x"04",
    x"10",x"00",x"40",x"00",x"80",x"09",x"00",x"0A",x"FF",x"33",x"00",x"00",x"05",x"50",x"16",x"0F",
    x"80",x"E1",x"02",x"80",x"00",x"07",x"04",x"54",x"AB",x"BE",x"AA",x"F5",x"BC",x"05",x"FF",x"00",
    x"07",x"EE",x"FF",x"BF",x"DF",x"EB",x"FF",x"E2",x"02",x"FD",x"00",x"01",x"F7",x"0E",x"FF",x"00",
    x"01",x"FE",x"05",x"FF",x"00",x"0F",x"EB",x"F7",x"C5",x"EF",x"EE",x"F8",x"FC",x"FF",x"0F",x"0B",
    x"1F",x"BE",x"F0",x"E0",x"80",x"4B",x"00",x"0A",x"FF",x"40",x"00",x"00",x"07",x"10",x"50",x"A0",
    x"F0",x"A8",x"F8",x"F0",x"06",x"F8",x"03",x"FC",x"00",x"04",x"FE",x"DC",x"FC",x"FE",x"04",x"FC",
    x"00",x"02",x"F8",x"F0",x"02",x"E0",x"02",x"80",x"00",x"02",x"00",x"80",x"03",x"00",x"00",x"01",
    x"80",x"03",x"C0",x"00",x"01",x"80",x"04",x"00",x"02",x"C0",x"00",x"01",x"80",x"38",x"00",x"00",
    x"01",x"01",x"16",x"00",x"0A",x"FF",x"45",x"00",x"02",x"03",x"00",x"02",x"05",x"03",x"05",x"07",
    x"00",x"02",x"0F",x"05",x"02",x"07",x"00",x"08",x"05",x"0E",x"0A",x"04",x"0B",x"15",x"05",x"01",
    x"05",x"00",x"00",x"03",x"01",x"07",x"01",x"46",x"00",x"00",x"01",x"02",x"15",x"00",x"0A",x"FF",
    x"31",x"00",x"00",x"08",x"05",x"07",x"1F",x"5F",x"2B",x"35",x"13",x"57",x"02",x"1F",x"00",x"02",
    x"FF",x"4F",x"02",x"05",x"00",x"07",x"07",x"5F",x"3F",x"5F",x"3F",x"1F",x"5F",x"0D",x"FF",x"00",
    x"02",x"7F",x"FF",x"02",x"7F",x"02",x"FF",x"00",x"05",x"1F",x"5F",x"17",x"1F",x"5F",x"02",x"7F",
    x"02",x"FF",x"00",x"03",x"7F",x"5F",x"7F",x"02",x"5F",x"00",x"02",x"0F",x"1F",x"02",x"17",x"00",
    x"04",x"15",x"07",x"00",x"01",x"3D",x"00",x"00",x"01",x"22",x"03",x"00",x"00",x"01",x"05",x"03",
    x"00",x"00",x"01",x"02",x"09",x"00",x"0A",x"FF",x"22",x"00",x"00",x"11",x"07",x"2F",x"7A",x"25",
    x"01",x"0B",x"07",x"0B",x"03",x"07",x"02",x"17",x"1F",x"3F",x"FF",x"AF",x"AB",x"33",x"FF",x"00",
    x"01",x"5F",x"06",x"FF",x"00",x"04",x"7F",x"5F",x"2F",x"0A",x"3E",x"00",x"02",x"40",x"02",x"54",
    x"02",x"55",x"00",x"03",x"5F",x"2A",x"AD",x"02",x"55",x"00",x"04",x"05",x"15",x"03",x"0A",x"0A",
    x"FF",x"1B",x"00",x"00",x"08",x"17",x"0A",x"17",x"28",x"7D",x"EB",x"F7",x"AB",x"0D",x"FF",x"00",
    x"01",x"BF",x"29",x"FF",x"00",x"01",x"FE",x"05",x"FF",x"00",x"01",x"FE",x"07",x"FF",x"00",x"01",
    x"FE",x"03",x"FF",x"00",x"0C",x"FE",x"FF",x"FE",x"FD",x"7D",x"BF",x"3F",x"3D",x"7B",x"55",x"2A",
    x"57",x"02",x"15",x"00",x"02",x"02",x"05",x"39",x"00",x"00",x"09",x"40",x"00",x"C0",x"40",x"E8",
    x"80",x"E8",x"54",x"5E",x"0A",x"FF",x"15",x"00",x"03",x"02",x"00",x"08",x"0B",x"0E",x"EF",x"FB",
    x"7F",x"2A",x"7F",x"AF",x"19",x"FF",x"00",x"16",x"FD",x"FE",x"F5",x"FF",x"D4",x"FE",x"FD",x"FA",
    x"F5",x"FA",x"D4",x"F6",x"AA",x"FA",x"A8",x"EA",x"D4",x"AC",x"A8",x"FA",x"F0",x"E8",x"02",x"E0",
    x"00",x"02",x"55",x"DF",x"04",x"FF",x"00",x"0E",x"F5",x"FF",x"55",x"FF",x"AB",x"7F",x"AF",x"FF",
    x"BD",x"D5",x"2A",x"55",x"A0",x"60",x"03",x"80",x"00",x"03",x"40",x"00",x"40",x"04",x"80",x"00",
    x"02",x"00",x"40",x"02",x"A0",x"00",x"19",x"00",x"A8",x"50",x"5A",x"AA",x"5E",x"A8",x"AD",x"04",
    x"55",x"42",x"5A",x"A8",x"2A",x"A8",x"AA",x"0A",x"56",x"AA",x"6A",x"A0",x"AA",x"05",x"AD",x"22",
    x"02",x"2A",x"00",x"04",x"0A",x"00",x"05",x"02",x"2C",x"00",x"0A",x"FF",x"0E",x"00",x"00",x"09",
    x"03",x"08",x"3D",x"15",x"55",x"2A",x"AF",x"AA",x"AF",x"02",x"FF",x"00",x"03",x"55",x"FF",x"AA",
    x"0F",x"FF",x"00",x"01",x"FD",x"05",x"FF",x"00",x"03",x"FD",x"FF",x"5F",x"05",x"FF",x"00",x"03",
    x"5F",x"D7",x"5F",x"02",x"54",x"00",x"07",x"24",x"00",x"40",x"00",x"80",x"00",x"80",x"0B",x"00",
    x"00",x"02",x"5A",x"FD",x"03",x"FF",x"00",x"05",x"7F",x"F7",x"A8",x"AA",x"F5",x"05",x"FF",x"02",
    x"AF",x"00",x"04",x"55",x"A5",x"14",x"15",x"11",x"00",x"00",x"03",x"AD",x"05",x"57",x"02",x"55",
    x"00",x"07",x"AA",x"AF",x"AA",x"BF",x"FD",x"F5",x"55",x"02",x"AF",x"00",x"01",x"FD",x"02",x"15",
    x"00",x"0F",x"05",x"C1",x"80",x"A0",x"80",x"F5",x"40",x"55",x"AA",x"AC",x"A8",x"B5",x"50",x"55",
    x"28",x"02",x"2A",x"00",x"02",x"0C",x"00",x"02",x"05",x"00",x"01",x"02",x"1A",x"00",x"00",x"07",
    x"01",x"03",x"00",x"07",x"00",x"0A",x"05",x"0A",x"FF",x"09",x"00",x"00",x"01",x"1F",x"03",x"00",
    x"00",x"05",x"5E",x"14",x"1A",x"AA",x"F5",x"02",x"FF",x"00",x"03",x"D5",x"FF",x"EF",x"05",x"FF",
    x"00",x"01",x"77",x"17",x"FF",x"00",x"04",x"FD",x"FE",x"E0",x"F0",x"02",x"80",x"17",x"00",x"05",
    x"FF",x"02",x"5F",x"00",x"01",x"57",x"03",x"FF",x"00",x"08",x"FB",x"FF",x"FD",x"FF",x"55",x"7B",
    x"54",x"F4",x"09",x"00",x"00",x"15",x"03",x"04",x"1A",x"14",x"A8",x"50",x"55",x"51",x"52",x"50",
    x"E0",x"80",x"F5",x"84",x"4A",x"55",x"6A",x"50",x"F5",x"75",x"7F",x"02",x"FF",x"00",x"19",x"7F",
    x"FF",x"BF",x"D7",x"55",x"5F",x"55",x"7A",x"13",x"57",x"04",x"57",x"15",x"7A",x"55",x"2A",x"00",
    x"55",x"04",x"6A",x"00",x"22",x"00",x"54",x"80",x"02",x"50",x"02",x"54",x"00",x"02",x"15",x"1D",
    x"02",x"15",x"00",x"05",x"07",x"05",x"07",x"02",x"07",x"03",x"05",x"00",x"10",x"15",x"0A",x"2A",
    x"17",x"3F",x"15",x"57",x"55",x"57",x"BF",x"AF",x"5F",x"BF",x"57",x"FF",x"3F",x"0B",x"FF",x"0A",
    x"00",x"00",x"0B",x"A0",x"28",x"10",x"14",x"00",x"0A",x"55",x"AF",x"15",x"BF",x"7F",x"1B",x"FF",
    x"00",x"04",x"EE",x"F5",x"40",x"80",x"1D",x"00",x"02",x"A0",x"00",x"03",x"F4",x"FA",x"FE",x"02",
    x"FF",x"00",x"03",x"BA",x"FF",x"EA",x"03",x"FF",x"00",x"05",x"FB",x"FF",x"EA",x"F8",x"40",x"10",
    x"00",x"02",x"0A",x"00",x"0C",x"57",x"3F",x"7F",x"15",x"AF",x"47",x"B5",x"0B",x"50",x"00",x"80",
    x"55",x"03",x"FF",x"00",x"16",x"AA",x"E8",x"54",x"FF",x"DF",x"FF",x"EB",x"EA",x"D4",x"A8",x"54",
    x"B5",x"02",x"D5",x"55",x"AA",x"55",x"AA",x"45",x"B5",x"00",x"A8",x"08",x"00",x"00",x"0F",x"40",
    x"EA",x"5B",x"AF",x"AA",x"FF",x"55",x"FF",x"57",x"FF",x"5F",x"FF",x"FD",x"FF",x"55",x"02",x"7F",
    x"03",x"FF",x"00",x"03",x"D5",x"FF",x"DF",x"03",x"FF",x"00",x"01",x"F5",x"0B",x"FF",x"0E",x"00",
    x"00",x"08",x"61",x"06",x"DF",x"AA",x"FF",x"55",x"FF",x"7F",x"18",x"FF",x"00",x"03",x"FE",x"AA",
    x"40",x"22",x"00",x"00",x"07",x"A0",x"40",x"80",x"40",x"80",x"C0",x"E0",x"03",x"C0",x"00",x"01",
    x"80",x"15",x"00",x"00",x"08",x"88",x"7A",x"54",x"F5",x"EA",x"7F",x"AA",x"7E",x"02",x"55",x"03",
    x"00",x"00",x"0B",x"FA",x"AA",x"FF",x"5B",x"C0",x"00",x"0A",x"80",x"FE",x"53",x"54",x"05",x"00",
    x"00",x"08",x"50",x"10",x"D7",x"FA",x"5F",x"AA",x"7A",x"55",x"0A",x"00",x"00",x"13",x"15",x"2A",
    x"AB",x"55",x"FF",x"AA",x"FF",x"FA",x"FF",x"55",x"FF",x"5F",x"BF",x"AA",x"F5",x"AA",x"FF",x"5F",
    x"EF",x"02",x"FF",x"00",x"07",x"AA",x"F7",x"5F",x"FF",x"7F",x"EF",x"EA",x"0A",x"FF",x"09",x"00",
    x"00",x"0D",x"01",x"06",x"54",x"5B",x"00",x"A0",x"2A",x"A5",x"5B",x"7F",x"EB",x"FA",x"EA",x"03",
    x"FF",x"00",x"01",x"FE",x"09",x"FF",x"00",x"01",x"FD",x"0B",x"FF",x"00",x"03",x"BF",x"2A",x"05",
    x"21",x"00",x"00",x"02",x"01",x"2F",x"02",x"55",x"00",x"04",x"0A",x"02",x"00",x"02",x"02",x"01",
    x"18",x"00",x"00",x"09",x"0A",x"0F",x"08",x"A0",x"40",x"6A",x"F8",x"E8",x"80",x"02",x"00",x"00",
    x"05",x"01",x"AA",x"EA",x"86",x"80",x"03",x"00",x"02",x"0A",x"00",x"01",x"A0",x"07",x"00",x"02",
    x"A0",x"00",x"04",x"FC",x"78",x"E8",x"80",x"0A",x"00",x"02",x"80",x"00",x"06",x"58",x"AA",x"FE",
    x"AA",x"FA",x"BE",x"03",x"FF",x"00",x"09",x"AA",x"FF",x"AA",x"FA",x"FF",x"D7",x"AA",x"D7",x"AA",
    x"02",x"7F",x"00",x"06",x"F5",x"AA",x"FF",x"AA",x"7F",x"5F",x"0A",x"FF",x"09",x"00",x"00",x"12",
    x"80",x"00",x"80",x"A8",x"57",x"AA",x"AF",x"AA",x"FF",x"BF",x"F7",x"FD",x"FF",x"AF",x"FF",x"BF",
    x"FF",x"DD",x"15",x"FF",x"00",x"03",x"0F",x"0B",x"02",x"1E",x"00",x"00",x"01",x"57",x"02",x"7F",
    x"02",x"FF",x"00",x"0C",x"55",x"FF",x"55",x"7F",x"5F",x"BF",x"AE",x"BF",x"55",x"57",x"15",x"05",
    x"0B",x"00",x"00",x"03",x"01",x"00",x"01",x"05",x"00",x"00",x"01",x"80",x"0A",x"00",x"00",x"04",
    x"A0",x"F7",x"45",x"02",x"03",x"00",x"00",x"02",x"85",x"88",x"1C",x"00",x"00",x"07",x"D5",x"54",
    x"EA",x"AA",x"EA",x"AA",x"BD",x"02",x"D5",x"02",x"AA",x"02",x"A8",x"00",x"0C",x"A4",x"BD",x"55",
    x"7A",x"A8",x"EA",x"F5",x"AA",x"F5",x"F7",x"A8",x"7A",x"0A",x"FF",x"0B",x"00",x"00",x"14",x"08",
    x"40",x"50",x"A0",x"5E",x"55",x"EA",x"45",x"EA",x"A8",x"FF",x"FD",x"FF",x"D5",x"FF",x"7F",x"FF",
    x"F5",x"FE",x"D5",x"09",x"FF",x"00",x"03",x"FB",x"FF",x"F7",x"07",x"FF",x"00",x"03",x"5F",x"FF",
    x"0B",x"02",x"02",x"19",x"00",x"00",x"02",x"03",x"BF",x"04",x"FF",x"00",x"03",x"FA",x"EC",x"FA",
    x"05",x"FF",x"00",x"06",x"7F",x"FA",x"00",x"D0",x"A0",x"56",x"0A",x"00",x"00",x"03",x"80",x"40",
    x"00",x"02",x"50",x"00",x"07",x"2A",x"54",x"28",x"0E",x"1F",x"05",x"0A",x"02",x"05",x"00",x"07",
    x"03",x"01",x"00",x"02",x"01",x"AA",x"FF",x"02",x"7F",x"00",x"03",x"FF",x"D1",x"02",x"1B",x"00",
    x"00",x"06",x"08",x"00",x"15",x"A0",x"56",x"00",x"02",x"50",x"00",x"0F",x"68",x"00",x"D0",x"00",
    x"40",x"00",x"40",x"00",x"A0",x"00",x"50",x"00",x"40",x"00",x"40",x"02",x"80",x"00",x"02",x"00",
    x"C0",x"0A",x"FF",x"0E",x"00",x"00",x"0C",x"04",x"17",x"AB",x"54",x"BC",x"54",x"D5",x"AA",x"EB",
    x"55",x"FF",x"7F",x"03",x"FF",x"00",x"03",x"5F",x"BF",x"7F",x"14",x"FF",x"00",x"09",x"BF",x"AB",
    x"D7",x"0F",x"57",x"07",x"0F",x"0B",x"05",x"12",x"00",x"00",x"06",x"14",x"F4",x"AA",x"F5",x"FC",
    x"FA",x"03",x"00",x"00",x"06",x"C0",x"AA",x"FF",x"5D",x"AF",x"08",x"1A",x"00",x"02",x"40",x"00",
    x"08",x"F0",x"40",x"50",x"E0",x"70",x"78",x"B8",x"70",x"02",x"F8",x"00",x"05",x"F0",x"50",x"A0",
    x"40",x"C0",x"2F",x"00",x"00",x"06",x"08",x"00",x"20",x"00",x"10",x"00",x"0A",x"FF",x"11",x"00",
    x"00",x"0D",x"07",x"08",x"80",x"C1",x"00",x"57",x"AA",x"7E",x"A8",x"EA",x"FB",x"FF",x"FA",x"0D",
    x"FF",x"00",x"01",x"AF",x"03",x"FF",x"00",x"02",x"D5",x"FF",x"02",x"FA",x"00",x"0B",x"E0",x"F0",
    x"E0",x"E8",x"D5",x"FD",x"E8",x"C0",x"FE",x"FF",x"85",x"14",x"00",x"00",x"01",x"50",x"08",x"00",
    x"00",x"03",x"80",x"40",x"80",x"60",x"00",x"0A",x"FF",x"11",x"00",x"00",x"02",x"70",x"02",x"02",
    x"A0",x"00",x"06",x"A8",x"A0",x"F5",x"D4",x"FA",x"AA",x"03",x"FF",x"00",x"01",x"F5",x"13",x"FF",
    x"00",x"11",x"57",x"FF",x"55",x"2F",x"BF",x"EF",x"5F",x"AF",x"15",x"D7",x"BF",x"FF",x"2E",x"0F",
    x"05",x"07",x"05",x"02",x"02",x"00",x"06",x"03",x"02",x"07",x"05",x"07",x"02",x"02",x"03",x"03",
    x"07",x"00",x"01",x"05",x"02",x"03",x"03",x"05",x"00",x"02",x"01",x"03",x"03",x"00",x"00",x"02",
    x"01",x"00",x"02",x"01",x"04",x"00",x"00",x"02",x"01",x"00",x"03",x"01",x"00",x"01",x"00",x"02",
    x"02",x"00",x"05",x"03",x"00",x"02",x"00",x"02",x"07",x"00",x"00",x"07",x"04",x"00",x"04",x"05",
    x"02",x"03",x"07",x"03",x"0F",x"00",x"04",x"1F",x"0F",x"1F",x"0F",x"02",x"1F",x"00",x"03",x"3F",
    x"7F",x"3F",x"02",x"3E",x"00",x"02",x"28",x"30",x"03",x"00",x"02",x"20",x"00",x"07",x"78",x"20",
    x"38",x"10",x"20",x"00",x"20",x"24",x"00",x"0A",x"FF",x"13",x"00",x"00",x"01",x"40",x"04",x"00",
    x"00",x"01",x"40",x"02",x"00",x"00",x"08",x"5C",x"54",x"7E",x"EB",x"EF",x"D5",x"FF",x"D5",x"11",
    x"FF",x"00",x"01",x"FA",x"09",x"FF",x"00",x"03",x"7F",x"FF",x"7F",x"03",x"FF",x"00",x"01",x"BF",
    x"17",x"FF",x"00",x"01",x"7F",x"07",x"FF",x"00",x"03",x"BF",x"FF",x"BF",x"06",x"FF",x"00",x"05",
    x"BF",x"AA",x"F5",x"20",x"1A",x"03",x"00",x"00",x"06",x"01",x"00",x"03",x"05",x"07",x"BE",x"02",
    x"FC",x"00",x"03",x"FE",x"F8",x"F0",x"04",x"F8",x"00",x"06",x"F0",x"F8",x"E0",x"F0",x"E8",x"F0",
    x"34",x"00",x"0A",x"FF",x"1E",x"00",x"00",x"0C",x"80",x"40",x"A0",x"E0",x"F4",x"54",x"F8",x"70",
    x"F8",x"EA",x"FF",x"EE",x"03",x"FF",x"00",x"07",x"FE",x"FD",x"EA",x"FD",x"F5",x"FF",x"DF",x"03",
    x"FF",x"00",x"02",x"FC",x"FE",x"03",x"FC",x"07",x"FF",x"00",x"01",x"DF",x"05",x"FF",x"00",x"01",
    x"D5",x"13",x"FF",x"00",x"03",x"F7",x"FF",x"D7",x"03",x"FF",x"00",x"01",x"FE",x"05",x"FF",x"00",
    x"01",x"AF",x"03",x"FF",x"00",x"09",x"F8",x"FC",x"50",x"7E",x"A8",x"F8",x"E0",x"EC",x"C0",x"03",
    x"80",x"45",x"00",x"0A",x"FF",x"2A",x"00",x"02",x"80",x"00",x"06",x"C0",x"80",x"22",x"6E",x"DC",
    x"08",x"04",x"00",x"00",x"0A",x"A0",x"40",x"50",x"28",x"10",x"20",x"E0",x"40",x"E0",x"CB",x"03",
    x"FF",x"00",x"02",x"FA",x"FE",x"02",x"FC",x"00",x"07",x"F3",x"FF",x"EA",x"FE",x"D4",x"F4",x"DC",
    x"02",x"FC",x"00",x"02",x"FE",x"EE",x"03",x"FF",x"00",x"05",x"FA",x"FE",x"F8",x"FE",x"F5",x"05",
    x"FF",x"00",x"02",x"F8",x"FC",x"02",x"F8",x"00",x"06",x"50",x"F4",x"54",x"F8",x"B8",x"F8",x"02",
    x"E0",x"02",x"C0",x"51",x"00",x"0A",x"FF",x"58",x"01",x"00",x"02",x"81",x"C1",x"02",x"81",x"62",
    x"01",x"C1",x"FF",x"08",x"00",x"00",x"00",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",
    x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",
    x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",
    x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",
    x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",
    x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",
    x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",
    x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",
    x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",
    x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",x"C8",x"C0",x"C7",x"08",
    x"C8",x"C0",x"C7",x"C8",x"C8",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"00",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"B7",x"A7",x"C0",x"B6",x"A7",x"C0",x"84",x"DF",x"20",
    x"F6",x"43",x"6F",x"75",x"63",x"6F",x"75",x"20",x"6C",x"65",x"73",x"20",x"70",x"69",x"72",x"61",
    x"74",x"65",x"73",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"00");

  CONSTANT ROM_BASIC6_2 : arr8 := (
    x"20",x"27",x"34",x"02",x"B6",x"A7",x"C0",x"84",x"DF",x"B7",x"A7",x"C0",x"35",x"02",x"AD",x"C4",
    x"34",x"02",x"B6",x"A7",x"C0",x"8A",x"20",x"B7",x"A7",x"C0",x"CE",x"DB",x"6D",x"34",x"40",x"20",
    x"EF",x"CE",x"DC",x"23",x"20",x"F7",x"32",x"62",x"39",x"CE",x"B0",x"A2",x"33",x"C5",x"EE",x"C5",
    x"C6",x"21",x"1F",x"9B",x"10",x"DF",x"75",x"AD",x"C4",x"5F",x"39",x"10",x"DE",x"75",x"39",x"BD",
    x"B0",x"8F",x"CC",x"B0",x"3B",x"DD",x"85",x"CC",x"D1",x"B3",x"FD",x"22",x"AE",x"0F",x"03",x"86",
    x"22",x"B7",x"20",x"1A",x"B7",x"20",x"1D",x"B7",x"20",x"1F",x"86",x"01",x"97",x"8A",x"CC",x"04",
    x"00",x"DD",x"9F",x"BD",x"E3",x"16",x"86",x"80",x"B7",x"22",x"B1",x"7D",x"20",x"80",x"27",x"03",
    x"BD",x"B2",x"4A",x"7E",x"DF",x"7F",x"CE",x"21",x"B7",x"20",x"A2",x"6E",x"9F",x"21",x"85",x"4D",
    x"27",x"1F",x"9B",x"8A",x"8D",x"03",x"90",x"8A",x"39",x"97",x"8B",x"B7",x"A7",x"E5",x"39",x"8E",
    x"22",x"B2",x"6F",x"82",x"8C",x"21",x"00",x"26",x"F9",x"86",x"06",x"97",x"8C",x"97",x"4D",x"97",
    x"30",x"39",x"B0",x"3F",x"B0",x"4D",x"B2",x"C8",x"B4",x"B7",x"B7",x"CE",x"B6",x"86",x"B6",x"E1",
    x"B8",x"FA",x"B3",x"AB",x"B3",x"A0",x"BC",x"88",x"BC",x"84",x"BB",x"89",x"BC",x"7E",x"B4",x"7F",
    x"B8",x"8D",x"B3",x"6A",x"B8",x"61",x"BA",x"F1",x"B8",x"B9",x"D3",x"FD",x"B4",x"16",x"DB",x"23",
    x"DE",x"A7",x"DF",x"96",x"E1",x"5B",x"E4",x"41",x"E7",x"56",x"E3",x"16",x"E7",x"B2",x"E2",x"34",
    x"E9",x"18",x"E9",x"1E",x"E9",x"2B",x"E9",x"37",x"E9",x"45",x"E9",x"4C",x"EA",x"2A",x"EA",x"62",
    x"EA",x"B0",x"EA",x"D5",x"C2",x"50",x"C3",x"01",x"C2",x"63",x"D1",x"B9",x"CF",x"9D",x"D0",x"55",
    x"CC",x"E2",x"CC",x"EB",x"CD",x"2D",x"CB",x"07",x"C2",x"F0",x"CA",x"B8",x"CC",x"44",x"CB",x"DD",
    x"CB",x"CF",x"CB",x"FF",x"CC",x"A9",x"C9",x"D6",x"CC",x"98",x"CC",x"6C",x"CC",x"B7",x"C1",x"84",
    x"C1",x"C4",x"C2",x"11",x"C4",x"0A",x"C5",x"18",x"C4",x"D4",x"CD",x"F0",x"EB",x"C1",x"EF",x"50",
    x"BC",x"AD",x"BB",x"90",x"B6",x"43",x"BD",x"B0",x"4D",x"7D",x"20",x"80",x"10",x"26",x"01",x"3A",
    x"39",x"BD",x"B0",x"3F",x"8E",x"23",x"00",x"6F",x"80",x"8C",x"2D",x"1F",x"23",x"F9",x"9F",x"1B",
    x"8E",x"9F",x"FF",x"9F",x"2E",x"8E",x"01",x"2C",x"9F",x"17",x"8E",x"2C",x"4E",x"BF",x"22",x"AE",
    x"B6",x"22",x"19",x"80",x"03",x"26",x"05",x"86",x"03",x"B7",x"2C",x"4D",x"B7",x"22",x"B0",x"8E",
    x"B0",x"76",x"9F",x"85",x"8E",x"2D",x"1D",x"9F",x"87",x"8E",x"23",x"2F",x"9F",x"97",x"8E",x"24",
    x"2F",x"9F",x"99",x"8E",x"B1",x"D6",x"8D",x"2F",x"8E",x"B2",x"05",x"8D",x"2A",x"8E",x"B1",x"C9",
    x"8D",x"25",x"8E",x"B8",x"F4",x"AF",x"43",x"AF",x"48",x"CE",x"27",x"A2",x"CC",x"7E",x"02",x"8D",
    x"1D",x"8E",x"BF",x"43",x"C6",x"0B",x"AF",x"C1",x"5A",x"26",x"FB",x"C6",x"02",x"8D",x"0F",x"CC",
    x"39",x"1B",x"8D",x"0A",x"8E",x"B1",x"F8",x"E6",x"1D",x"EE",x"1E",x"7E",x"DF",x"87",x"A7",x"C0",
    x"AF",x"C1",x"5A",x"26",x"F9",x"39",x"0A",x"27",x"70",x"79",x"D8",x"0C",x"B0",x"E5",x"41",x"D9",
    x"F1",x"B0",x"3D",x"1F",x"21",x"B7",x"7E",x"B2",x"07",x"7E",x"B8",x"DD",x"7E",x"B8",x"DF",x"0C",
    x"C8",x"26",x"02",x"0C",x"C7",x"B6",x"00",x"00",x"81",x"20",x"27",x"F3",x"81",x"3A",x"24",x"04",
    x"80",x"30",x"80",x"D0",x"39",x"0A",x"29",x"1A",x"DC",x"AB",x"DC",x"CC",x"DE",x"99",x"DD",x"5C",
    x"DE",x"19",x"2F",x"23",x"00",x"C6",x"05",x"27",x"1B",x"7A",x"23",x"01",x"26",x"25",x"F6",x"2B",
    x"3B",x"27",x"11",x"8E",x"00",x"00",x"27",x"0C",x"30",x"1F",x"BF",x"23",x"0F",x"26",x"05",x"C6",
    x"FF",x"F7",x"2B",x"34",x"8E",x"00",x"00",x"27",x"0A",x"30",x"1F",x"BF",x"23",x"20",x"26",x"03",
    x"73",x"22",x"A9",x"3B",x"28",x"50",x"11",x"80",x"28",x"50",x"11",x"FF",x"50",x"A0",x"11",x"FF",
    x"19",x"32",x"FF",x"80",x"9C",x"A1",x"C6",x"D3",x"EA",x"C3",x"8E",x"B2",x"44",x"C6",x"07",x"86",
    x"02",x"5A",x"2B",x"0B",x"B6",x"A0",x"03",x"48",x"48",x"A8",x"85",x"85",x"FC",x"26",x"F0",x"B7",
    x"22",x"19",x"C6",x"04",x"3D",x"8E",x"B2",x"34",x"3A",x"EC",x"81",x"FD",x"22",x"1F",x"EC",x"84",
    x"B7",x"22",x"23",x"F7",x"22",x"B1",x"C6",x"01",x"20",x"40",x"CC",x"03",x"07",x"B1",x"22",x"19",
    x"27",x"01",x"5F",x"F7",x"20",x"4B",x"4F",x"B7",x"20",x"49",x"4C",x"B7",x"20",x"4C",x"9E",x"97",
    x"BF",x"20",x"4F",x"8D",x"23",x"24",x"1D",x"B6",x"20",x"4E",x"84",x"8E",x"27",x"15",x"BD",x"B3",
    x"8B",x"27",x"10",x"C6",x"04",x"8D",x"13",x"8D",x"0F",x"25",x"06",x"C6",x"80",x"F7",x"22",x"B1",
    x"39",x"8D",x"02",x"43",x"39",x"C6",x"10",x"8C",x"C6",x"02",x"F7",x"20",x"48",x"3F",x"A6",x"BF",
    x"27",x"6D",x"1F",x"98",x"10",x"8E",x"00",x"05",x"4A",x"97",x"95",x"CE",x"22",x"24",x"AF",x"C1",
    x"6F",x"84",x"30",x"89",x"01",x"1B",x"4A",x"2A",x"F5",x"9E",x"99",x"CC",x"00",x"A6",x"6F",x"84",
    x"30",x"8B",x"31",x"3F",x"26",x"F8",x"39",x"0C",x"89",x"8D",x"15",x"7E",x"EF",x"81",x"B7",x"20",
    x"4B",x"F7",x"20",x"4C",x"C6",x"08",x"20",x"08",x"B7",x"20",x"4B",x"F7",x"20",x"4C",x"C6",x"02",
    x"9E",x"97",x"BF",x"20",x"4F",x"F7",x"20",x"48",x"7E",x"ED",x"D3",x"8E",x"B3",x"19",x"B6",x"20",
    x"4E",x"E6",x"80",x"44",x"24",x"FB",x"7E",x"BD",x"91",x"48",x"35",x"35",x"35",x"47",x"4B",x"35",
    x"4C",x"34",x"16",x"8D",x"2E",x"6F",x"01",x"30",x"05",x"6F",x"84",x"C6",x"08",x"8D",x"D3",x"35",
    x"96",x"8D",x"20",x"6D",x"84",x"27",x"01",x"39",x"6F",x"01",x"33",x"05",x"8D",x"C0",x"30",x"01",
    x"F6",x"22",x"20",x"3A",x"86",x"FE",x"8C",x"A7",x"80",x"5C",x"26",x"FB",x"9E",x"97",x"C6",x"A1",
    x"7E",x"DF",x"87",x"CC",x"14",x"02",x"B7",x"20",x"4B",x"F7",x"20",x"4C",x"34",x"06",x"B6",x"20",
    x"49",x"C6",x"A6",x"3D",x"9E",x"99",x"30",x"8B",x"35",x"86",x"8D",x"C5",x"8D",x"EE",x"30",x"06",
    x"6F",x"E2",x"C6",x"A0",x"A6",x"80",x"43",x"26",x"02",x"6C",x"E4",x"5A",x"26",x"F6",x"4F",x"8D",
    x"0A",x"27",x"03",x"68",x"E4",x"49",x"35",x"04",x"7E",x"CB",x"03",x"F6",x"22",x"B1",x"C1",x"80",
    x"39",x"0F",x"8E",x"86",x"14",x"B7",x"20",x"4B",x"8D",x"F1",x"4F",x"D3",x"97",x"DD",x"F1",x"39",
    x"96",x"8E",x"B7",x"20",x"4C",x"8D",x"EA",x"9E",x"8F",x"20",x"46",x"17",x"FF",x"83",x"0F",x"92",
    x"9E",x"97",x"9F",x"8F",x"8D",x"DB",x"C6",x"03",x"BD",x"B2",x"FB",x"9F",x"8F",x"A6",x"84",x"27",
    x"2E",x"43",x"27",x"1F",x"CE",x"22",x"4F",x"C6",x"0A",x"A6",x"C5",x"27",x"04",x"A1",x"85",x"26",
    x"20",x"5A",x"2A",x"F5",x"B6",x"20",x"4C",x"97",x"8E",x"E6",x"0D",x"D7",x"91",x"8D",x"22",x"34",
    x"02",x"20",x"9B",x"D6",x"92",x"26",x"07",x"F6",x"20",x"4C",x"D7",x"92",x"9F",x"93",x"39",x"8D",
    x"F2",x"30",x"88",x"20",x"9C",x"F1",x"25",x"C3",x"F6",x"20",x"4C",x"5C",x"C1",x"10",x"23",x"B8",
    x"39",x"BD",x"B3",x"5C",x"33",x"06",x"4F",x"4C",x"10",x"27",x"01",x"9A",x"1F",x"31",x"3A",x"E6",
    x"84",x"C1",x"C0",x"25",x"F2",x"39",x"CC",x"14",x"01",x"BD",x"B2",x"F8",x"C6",x"08",x"D7",x"51",
    x"6D",x"84",x"2A",x"F1",x"33",x"84",x"8E",x"B4",x"2C",x"7E",x"DF",x"87",x"4E",x"6F",x"20",x"4E",
    x"61",x"6D",x"65",x"20",x"34",x"02",x"D6",x"95",x"8D",x"2A",x"27",x"15",x"B6",x"20",x"49",x"A1",
    x"01",x"26",x"0E",x"DE",x"8F",x"A6",x"4D",x"A1",x"02",x"26",x"06",x"A6",x"84",x"A1",x"E4",x"27",
    x"29",x"5A",x"2A",x"E4",x"35",x"82",x"BD",x"B3",x"AB",x"0D",x"8E",x"26",x"1A",x"39",x"34",x"04",
    x"F6",x"22",x"44",x"8C",x"34",x"04",x"58",x"8E",x"22",x"24",x"AE",x"85",x"E6",x"84",x"35",x"84",
    x"0D",x"8E",x"26",x"E9",x"C6",x"3E",x"8C",x"C6",x"42",x"8C",x"C6",x"34",x"7E",x"BD",x"91",x"0C",
    x"89",x"BD",x"B3",x"AB",x"8D",x"EA",x"8D",x"03",x"7E",x"EF",x"81",x"86",x"FF",x"8D",x"A5",x"6F",
    x"9F",x"21",x"8F",x"BD",x"B2",x"F4",x"D6",x"91",x"BD",x"B3",x"5C",x"33",x"06",x"86",x"FF",x"1F",
    x"31",x"3A",x"E6",x"84",x"A7",x"84",x"C1",x"C0",x"25",x"F5",x"7E",x"B3",x"21",x"0C",x"89",x"D6",
    x"95",x"96",x"77",x"81",x"11",x"26",x"06",x"D6",x"95",x"8D",x"A9",x"27",x"08",x"5A",x"2A",x"F9",
    x"C6",x"40",x"7E",x"BD",x"91",x"F7",x"22",x"44",x"BF",x"22",x"45",x"BD",x"B3",x"AB",x"B6",x"22",
    x"4B",x"81",x"20",x"26",x"13",x"96",x"8E",x"27",x"08",x"97",x"92",x"9E",x"8F",x"9F",x"93",x"8D",
    x"AA",x"BD",x"B5",x"F6",x"8D",x"59",x"20",x"1F",x"81",x"10",x"26",x"29",x"8D",x"82",x"BD",x"B4",
    x"34",x"9E",x"8F",x"EC",x"0B",x"FD",x"22",x"4C",x"30",x"88",x"10",x"CE",x"22",x"91",x"C6",x"10",
    x"BD",x"DF",x"87",x"8D",x"30",x"8D",x"6C",x"BD",x"B3",x"5C",x"6C",x"84",x"BE",x"22",x"45",x"B6",
    x"22",x"4B",x"A7",x"84",x"39",x"96",x"8E",x"26",x"05",x"BD",x"B5",x"F6",x"20",x"05",x"86",x"FF",
    x"BD",x"B4",x"34",x"8D",x"10",x"63",x"0D",x"6C",x"08",x"FE",x"22",x"AA",x"EF",x"0B",x"FC",x"22",
    x"47",x"ED",x"09",x"20",x"D2",x"8D",x"08",x"DE",x"8F",x"EE",x"4E",x"EF",x"88",x"13",x"39",x"BE",
    x"22",x"45",x"C6",x"1B",x"6F",x"80",x"5A",x"26",x"FB",x"BE",x"22",x"45",x"BD",x"B3",x"8B",x"E7",
    x"88",x"1A",x"B6",x"20",x"49",x"A7",x"01",x"96",x"91",x"A7",x"02",x"A7",x"03",x"D6",x"8E",x"C0",
    x"03",x"58",x"58",x"58",x"34",x"04",x"DC",x"8F",x"93",x"97",x"86",x"08",x"3D",x"AB",x"E0",x"A7",
    x"88",x"12",x"39",x"6F",x"05",x"A6",x"01",x"B7",x"20",x"49",x"A6",x"04",x"4C",x"34",x"02",x"81",
    x"08",x"23",x"01",x"4F",x"A7",x"04",x"E6",x"03",x"33",x"84",x"BD",x"B3",x"5C",x"3A",x"E6",x"06",
    x"30",x"C4",x"C1",x"C0",x"24",x"0A",x"35",x"02",x"80",x"09",x"26",x"15",x"E7",x"03",x"20",x"DC",
    x"C4",x"3F",x"C1",x"08",x"23",x"05",x"C6",x"46",x"7E",x"BD",x"91",x"E0",x"E0",x"25",x"14",x"1F",
    x"98",x"34",x"02",x"8D",x"16",x"8D",x"2C",x"E6",x"88",x"1A",x"6D",x"E0",x"26",x"09",x"EC",x"88",
    x"13",x"26",x"04",x"5F",x"63",x"88",x"17",x"E7",x"88",x"18",x"39",x"6C",x"08",x"26",x"02",x"6C",
    x"07",x"39",x"E6",x"03",x"86",x"08",x"54",x"F7",x"20",x"4B",x"25",x"01",x"4F",x"AB",x"04",x"B7",
    x"20",x"4C",x"39",x"C6",x"02",x"8C",x"C6",x"08",x"F7",x"20",x"48",x"8D",x"E5",x"33",x"88",x"1B",
    x"FF",x"20",x"4F",x"7E",x"ED",x"D3",x"D6",x"92",x"26",x"05",x"C6",x"41",x"7E",x"BD",x"91",x"D7",
    x"8E",x"BD",x"B2",x"FB",x"9E",x"93",x"9F",x"8F",x"33",x"84",x"C6",x"20",x"6F",x"80",x"5A",x"26",
    x"FB",x"34",x"40",x"BD",x"B8",x"7E",x"33",x"45",x"C6",x"08",x"BD",x"DF",x"87",x"35",x"40",x"FC",
    x"22",x"4C",x"ED",x"4B",x"C6",x"27",x"BD",x"B7",x"81",x"97",x"91",x"A7",x"4D",x"BD",x"B2",x"F4",
    x"34",x"76",x"BD",x"B3",x"5C",x"6C",x"01",x"A6",x"01",x"B1",x"22",x"23",x"25",x"03",x"BD",x"B3",
    x"21",x"35",x"F6",x"0F",x"78",x"9F",x"50",x"BD",x"B4",x"5E",x"E6",x"88",x"17",x"26",x"70",x"E6",
    x"05",x"4F",x"33",x"8B",x"33",x"C8",x"1B",x"E6",x"88",x"18",x"34",x"10",x"9E",x"50",x"27",x"0B",
    x"A6",x"C0",x"A7",x"A0",x"5A",x"27",x"14",x"30",x"1F",x"26",x"F5",x"9F",x"50",x"AE",x"E4",x"E7",
    x"88",x"18",x"1F",x"30",x"A3",x"E1",x"C0",x"1B",x"E7",x"05",x"39",x"30",x"1F",x"9F",x"50",x"35",
    x"10",x"BD",x"B5",x"73",x"20",x"C4",x"0F",x"78",x"F6",x"22",x"44",x"58",x"8E",x"22",x"24",x"AE",
    x"85",x"E6",x"84",x"C1",x"40",x"26",x"16",x"EC",x"88",x"15",x"10",x"A3",x"09",x"24",x"20",x"C3",
    x"00",x"01",x"ED",x"88",x"15",x"AE",x"0B",x"30",x"8B",x"A6",x"1F",x"20",x"22",x"E6",x"88",x"10",
    x"27",x"08",x"A6",x"88",x"11",x"6F",x"88",x"10",x"20",x"15",x"E6",x"88",x"17",x"27",x"03",x"03",
    x"78",x"39",x"E6",x"05",x"6C",x"05",x"6A",x"88",x"18",x"27",x"07",x"3A",x"A6",x"88",x"1B",x"97",
    x"96",x"39",x"4F",x"33",x"8B",x"A6",x"C8",x"1B",x"97",x"96",x"34",x"02",x"BD",x"B5",x"73",x"35",
    x"82",x"BD",x"B4",x"5E",x"BF",x"22",x"45",x"A6",x"84",x"27",x"E6",x"34",x"02",x"6F",x"84",x"E6",
    x"01",x"F7",x"20",x"49",x"81",x"10",x"27",x"1F",x"81",x"20",x"26",x"1B",x"E6",x"88",x"18",x"86",
    x"80",x"6D",x"05",x"27",x"03",x"E6",x"88",x"1A",x"ED",x"88",x"13",x"6C",x"04",x"E6",x"03",x"BD",
    x"B3",x"5C",x"A7",x"01",x"3A",x"6C",x"06",x"BD",x"B3",x"5C",x"6A",x"84",x"6D",x"01",x"27",x"03",
    x"BD",x"B3",x"21",x"BE",x"22",x"45",x"35",x"02",x"81",x"20",x"27",x"08",x"81",x"40",x"26",x"06",
    x"A6",x"0F",x"27",x"08",x"8D",x"03",x"7E",x"EF",x"81",x"BD",x"B5",x"E6",x"A6",x"88",x"13",x"2A",
    x"90",x"E6",x"88",x"12",x"C4",x"07",x"86",x"20",x"3D",x"DE",x"97",x"31",x"CB",x"E6",x"88",x"12",
    x"54",x"54",x"54",x"CB",x"03",x"86",x"14",x"BD",x"B2",x"F8",x"BE",x"22",x"45",x"EC",x"88",x"13",
    x"84",x"7F",x"ED",x"2E",x"7D",x"22",x"4A",x"27",x"15",x"C6",x"10",x"8E",x"22",x"91",x"33",x"A8",
    x"10",x"6D",x"C4",x"27",x"06",x"30",x"08",x"33",x"48",x"C0",x"08",x"BD",x"DF",x"87",x"7E",x"B2",
    x"F4",x"34",x"40",x"BD",x"B3",x"5C",x"33",x"06",x"4F",x"C4",x"FE",x"6F",x"E2",x"30",x"C4",x"3A",
    x"63",x"84",x"27",x"30",x"63",x"84",x"4C",x"81",x"A0",x"24",x"25",x"5C",x"C5",x"01",x"26",x"ED",
    x"34",x"06",x"C0",x"02",x"63",x"62",x"26",x"0C",x"E0",x"E0",x"2A",x"04",x"E6",x"E4",x"63",x"61",
    x"32",x"61",x"20",x"D9",x"EB",x"E0",x"C1",x"A0",x"25",x"F6",x"E6",x"E4",x"C0",x"04",x"20",x"EE",
    x"C6",x"3F",x"20",x"38",x"32",x"61",x"1F",x"98",x"C6",x"C0",x"E7",x"84",x"35",x"C0",x"F6",x"22",
    x"44",x"58",x"8E",x"22",x"24",x"AE",x"85",x"E6",x"84",x"C1",x"10",x"27",x"2D",x"81",x"0D",x"26",
    x"02",x"6F",x"06",x"81",x"20",x"25",x"02",x"6C",x"06",x"C1",x"40",x"26",x"1E",x"34",x"02",x"EC",
    x"88",x"17",x"C3",x"00",x"01",x"10",x"A3",x"09",x"23",x"05",x"C6",x"4A",x"7E",x"BD",x"91",x"ED",
    x"88",x"17",x"AE",x"0B",x"30",x"8B",x"35",x"02",x"A7",x"1F",x"39",x"6C",x"88",x"18",x"E6",x"88",
    x"18",x"34",x"10",x"3A",x"A7",x"88",x"1A",x"35",x"10",x"E1",x"88",x"1A",x"27",x"01",x"39",x"6F",
    x"88",x"18",x"E6",x"01",x"F7",x"20",x"49",x"6C",x"04",x"BD",x"B7",x"39",x"31",x"84",x"E6",x"03",
    x"BD",x"B3",x"5C",x"3A",x"33",x"06",x"A6",x"24",x"81",x"08",x"25",x"0E",x"6A",x"24",x"6C",x"25",
    x"BD",x"B7",x"81",x"6F",x"24",x"6F",x"25",x"A7",x"23",x"8C",x"8A",x"C0",x"A7",x"C4",x"30",x"A4",
    x"BD",x"B5",x"CB",x"7E",x"B6",x"30",x"BD",x"B4",x"64",x"A6",x"06",x"5F",x"1F",x"01",x"86",x"0E",
    x"39",x"BD",x"EF",x"67",x"DE",x"97",x"FF",x"20",x"4F",x"96",x"8D",x"B7",x"20",x"48",x"3F",x"2A",
    x"10",x"25",x"FA",x"97",x"8D",x"08",x"CC",x"14",x"01",x"BD",x"B2",x"EE",x"20",x"35",x"8E",x"22",
    x"4F",x"C6",x"0B",x"20",x"05",x"CE",x"22",x"4F",x"C6",x"13",x"7E",x"DF",x"87",x"34",x"30",x"1F",
    x"21",x"8D",x"F2",x"BD",x"B4",x"56",x"35",x"10",x"8D",x"EB",x"BD",x"B3",x"AB",x"BD",x"B4",x"70",
    x"35",x"10",x"DE",x"8F",x"8D",x"DB",x"33",x"45",x"6D",x"84",x"27",x"04",x"C6",x"08",x"8D",x"DA",
    x"BD",x"B2",x"F4",x"7E",x"EF",x"81",x"F6",x"22",x"44",x"BD",x"B4",x"64",x"EC",x"07",x"7E",x"CB",
    x"03",x"F6",x"22",x"44",x"BD",x"B4",x"64",x"CC",x"10",x"33",x"A1",x"84",x"10",x"26",x"04",x"C1",
    x"5F",x"A6",x"88",x"10",x"26",x"03",x"E6",x"88",x"17",x"7E",x"C2",x"52",x"34",x"14",x"BD",x"B4",
    x"5E",x"E6",x"84",x"C1",x"40",x"26",x"0B",x"EC",x"88",x"15",x"83",x"00",x"01",x"ED",x"88",x"15",
    x"35",x"94",x"A7",x"88",x"11",x"63",x"88",x"10",x"35",x"94",x"34",x"10",x"BD",x"B4",x"5E",x"BF",
    x"22",x"45",x"6F",x"88",x"15",x"6F",x"88",x"16",x"6F",x"88",x"17",x"6F",x"88",x"18",x"6F",x"06",
    x"A6",x"01",x"B7",x"20",x"49",x"EC",x"E1",x"27",x"02",x"ED",x"07",x"EE",x"07",x"BD",x"B5",x"CB",
    x"EC",x"09",x"AE",x"0B",x"34",x"16",x"30",x"5F",x"BD",x"BA",x"BD",x"34",x"60",x"A6",x"E0",x"26",
    x"1E",x"BD",x"B3",x"8B",x"26",x"10",x"68",x"62",x"69",x"61",x"69",x"E4",x"25",x"11",x"64",x"62",
    x"35",x"10",x"35",x"04",x"20",x"04",x"35",x"12",x"8D",x"0A",x"8C",x"05",x"00",x"25",x"2F",x"C6",
    x"45",x"7E",x"BD",x"91",x"34",x"12",x"AE",x"E4",x"E6",x"62",x"3A",x"34",x"10",x"1F",x"10",x"EB",
    x"E4",x"24",x"08",x"CB",x"01",x"AE",x"62",x"30",x"01",x"AF",x"62",x"E7",x"61",x"AE",x"62",x"E6",
    x"E0",x"3A",x"E6",x"E0",x"53",x"26",x"03",x"30",x"01",x"86",x"53",x"32",x"63",x"39",x"FE",x"22",
    x"45",x"AC",x"4D",x"10",x"27",x"00",x"A6",x"34",x"14",x"A6",x"4F",x"27",x"06",x"6F",x"4F",x"C6",
    x"08",x"8D",x"34",x"EC",x"61",x"BD",x"BA",x"E7",x"34",x"04",x"17",x"01",x"19",x"50",x"EB",x"63",
    x"5C",x"E7",x"44",x"E6",x"42",x"BD",x"B3",x"5C",x"33",x"06",x"A6",x"E4",x"4C",x"30",x"C4",x"3A",
    x"4A",x"27",x"36",x"E7",x"E4",x"E6",x"84",x"C1",x"C0",x"25",x"F2",x"E6",x"E4",x"7D",x"22",x"49",
    x"26",x"16",x"C6",x"36",x"7E",x"BD",x"91",x"30",x"C8",x"1B",x"F7",x"20",x"48",x"BF",x"20",x"4F",
    x"30",x"C4",x"BD",x"B5",x"D2",x"7E",x"ED",x"D3",x"34",x"12",x"BD",x"B7",x"81",x"1F",x"89",x"35",
    x"42",x"E7",x"C4",x"4A",x"26",x"F2",x"BD",x"B3",x"21",x"32",x"61",x"FE",x"22",x"45",x"E7",x"43",
    x"86",x"FF",x"A7",x"4D",x"A6",x"84",x"81",x"C0",x"25",x"2B",x"84",x"3F",x"A1",x"44",x"24",x"25",
    x"B6",x"22",x"49",x"27",x"BD",x"A6",x"44",x"8A",x"C0",x"A7",x"84",x"BD",x"B6",x"30",x"AE",x"63",
    x"AC",x"C8",x"19",x"26",x"0B",x"AC",x"C8",x"13",x"27",x"0B",x"E6",x"C8",x"1A",x"86",x"80",x"8C",
    x"4F",x"5F",x"ED",x"C8",x"13",x"C6",x"02",x"8D",x"9E",x"35",x"14",x"AF",x"4D",x"34",x"04",x"BD",
    x"B3",x"5C",x"30",x"06",x"E6",x"43",x"3A",x"A6",x"84",x"81",x"C0",x"25",x"2D",x"84",x"3F",x"A1",
    x"44",x"26",x"27",x"EC",x"C8",x"13",x"84",x"7F",x"34",x"06",x"4F",x"E6",x"62",x"E3",x"63",x"10",
    x"A3",x"E1",x"23",x"16",x"7D",x"22",x"49",x"10",x"27",x"FF",x"67",x"1F",x"01",x"AC",x"C8",x"19",
    x"23",x"03",x"EC",x"C8",x"19",x"8A",x"80",x"ED",x"C8",x"13",x"35",x"04",x"30",x"C8",x"1B",x"3A",
    x"34",x"04",x"E6",x"C8",x"1A",x"E0",x"E4",x"86",x"FF",x"50",x"E3",x"61",x"24",x"09",x"ED",x"61",
    x"E6",x"C8",x"1A",x"E0",x"E0",x"20",x"08",x"E6",x"62",x"6F",x"61",x"6F",x"62",x"32",x"61",x"EE",
    x"62",x"B6",x"22",x"49",x"27",x"02",x"1E",x"13",x"BD",x"DF",x"87",x"EF",x"62",x"FE",x"22",x"45",
    x"B6",x"22",x"49",x"27",x"04",x"A7",x"4F",x"AF",x"62",x"AE",x"4D",x"30",x"01",x"5F",x"EE",x"E4",
    x"10",x"26",x"FE",x"96",x"35",x"96",x"58",x"49",x"58",x"49",x"58",x"49",x"39",x"34",x"76",x"6F",
    x"64",x"A6",x"63",x"3D",x"ED",x"66",x"EC",x"61",x"3D",x"EB",x"66",x"89",x"00",x"ED",x"65",x"E6",
    x"E4",x"A6",x"63",x"3D",x"E3",x"65",x"ED",x"65",x"24",x"02",x"6C",x"64",x"A6",x"E4",x"E6",x"62",
    x"3D",x"E3",x"64",x"ED",x"64",x"35",x"F6",x"44",x"56",x"44",x"56",x"44",x"56",x"39",x"F7",x"22",
    x"44",x"BD",x"B4",x"5E",x"A6",x"01",x"B7",x"20",x"49",x"E6",x"02",x"34",x"10",x"BD",x"B4",x"01",
    x"4A",x"C4",x"3F",x"34",x"04",x"1F",x"89",x"4F",x"8D",x"AC",x"EB",x"E0",x"89",x"00",x"35",x"10",
    x"34",x"02",x"A6",x"84",x"81",x"40",x"35",x"02",x"10",x"26",x"0F",x"E7",x"34",x"10",x"83",x"00",
    x"00",x"27",x"03",x"83",x"00",x"01",x"8D",x"31",x"8E",x"BD",x"EE",x"BD",x"B3",x"8B",x"26",x"02",
    x"30",x"04",x"BD",x"BF",x"6A",x"BD",x"C2",x"11",x"AE",x"E4",x"EC",x"88",x"13",x"84",x"7F",x"8D",
    x"18",x"8E",x"BE",x"0B",x"BD",x"CB",x"C1",x"BD",x"C2",x"11",x"35",x"10",x"EC",x"09",x"8D",x"09",
    x"8E",x"C0",x"BB",x"BD",x"CB",x"C1",x"7E",x"C3",x"01",x"1F",x"01",x"7E",x"CB",x"91",x"34",x"12",
    x"9E",x"1F",x"96",x"21",x"30",x"01",x"9F",x"6B",x"97",x"6D",x"9E",x"25",x"96",x"27",x"9F",x"6E",
    x"97",x"70",x"35",x"92",x"D3",x"6B",x"93",x"6E",x"24",x"01",x"39",x"C6",x"07",x"7E",x"BD",x"91",
    x"BD",x"B8",x"85",x"E6",x"84",x"F7",x"20",x"49",x"39",x"0F",x"6D",x"0F",x"70",x"8C",x"8D",x"CE",
    x"B6",x"22",x"B0",x"97",x"FD",x"CC",x"FF",x"FF",x"DD",x"F6",x"B7",x"22",x"4A",x"0F",x"9D",x"10",
    x"9F",x"FB",x"9C",x"FB",x"26",x"02",x"03",x"9D",x"8D",x"D6",x"86",x"10",x"97",x"F8",x"17",x"00",
    x"B0",x"D7",x"F6",x"9E",x"50",x"9F",x"F9",x"BD",x"EF",x"B5",x"D6",x"F6",x"F7",x"22",x"44",x"9E",
    x"6E",x"96",x"70",x"9F",x"F3",x"97",x"F5",x"8D",x"73",x"8D",x"7D",x"24",x"11",x"34",x"14",x"BD",
    x"B6",x"86",x"35",x"14",x"0D",x"78",x"26",x"04",x"A7",x"80",x"20",x"ED",x"8D",x"7C",x"9F",x"F3",
    x"D7",x"F5",x"0D",x"9D",x"27",x"03",x"17",x"00",x"85",x"0D",x"F8",x"27",x"1A",x"9E",x"FB",x"8D",
    x"8F",x"BD",x"B3",x"6A",x"DC",x"50",x"93",x"F9",x"10",x"25",x"FB",x"C4",x"BD",x"B4",x"56",x"86",
    x"20",x"8D",x"5E",x"D7",x"F7",x"0F",x"F8",x"BD",x"EF",x"B5",x"D6",x"F7",x"F7",x"22",x"44",x"8D",
    x"2B",x"8D",x"35",x"24",x"0B",x"A6",x"80",x"34",x"14",x"BD",x"B7",x"CE",x"35",x"14",x"20",x"F1",
    x"D6",x"78",x"26",x"0B",x"0D",x"9D",x"27",x"05",x"BD",x"B3",x"21",x"8D",x"41",x"20",x"88",x"96",
    x"FD",x"B7",x"22",x"B0",x"8D",x"24",x"7F",x"22",x"4A",x"0F",x"9D",x"39",x"9E",x"6B",x"D6",x"6D",
    x"1E",x"98",x"BD",x"B0",x"7F",x"1E",x"98",x"39",x"8C",x"9E",x"FF",x"23",x"06",x"8E",x"60",x"00",
    x"5C",x"8D",x"ED",x"D1",x"F5",x"26",x"02",x"9C",x"F3",x"39",x"34",x"76",x"BD",x"B6",x"E1",x"35",
    x"F6",x"34",x"72",x"B7",x"22",x"4B",x"BD",x"B4",x"B7",x"F6",x"22",x"44",x"35",x"F2",x"BD",x"EF",
    x"81",x"BD",x"EF",x"67",x"96",x"FD",x"B7",x"22",x"B0",x"35",x"10",x"9F",x"9B",x"39",x"BD",x"B3",
    x"53",x"BD",x"B3",x"38",x"6E",x"9F",x"21",x"9B",x"B1",x"20",x"49",x"27",x"06",x"0F",x"6D",x"0F",
    x"70",x"20",x"1A",x"8E",x"60",x"00",x"86",x"01",x"9F",x"6B",x"97",x"6D",x"8E",x"9F",x"FF",x"96",
    x"8C",x"9F",x"6E",x"97",x"70",x"B6",x"20",x"49",x"20",x"03",x"BD",x"BB",x"5E",x"F6",x"20",x"49",
    x"DD",x"8E",x"4F",x"BD",x"B3",x"8B",x"27",x"02",x"5F",x"4C",x"DD",x"90",x"0F",x"9D",x"96",x"8E",
    x"91",x"8F",x"26",x"02",x"03",x"9D",x"CC",x"00",x"01",x"DD",x"92",x"9E",x"6E",x"96",x"70",x"30",
    x"89",x"FF",x"00",x"8C",x"60",x"00",x"24",x"04",x"8E",x"9E",x"FF",x"4A",x"9F",x"F3",x"97",x"F5",
    x"96",x"8E",x"B7",x"20",x"49",x"86",x"02",x"B7",x"20",x"48",x"8D",x"2E",x"9F",x"F3",x"D7",x"F5",
    x"0D",x"9D",x"27",x"02",x"8D",x"83",x"96",x"8F",x"B7",x"20",x"49",x"86",x"08",x"B7",x"20",x"48",
    x"8D",x"18",x"B6",x"20",x"4B",x"F6",x"20",x"4C",x"DD",x"92",x"0D",x"78",x"26",x"09",x"0D",x"9D",
    x"27",x"03",x"BD",x"BC",x"79",x"20",x"B4",x"0F",x"9D",x"39",x"BD",x"EE",x"51",x"0F",x"78",x"DC",
    x"92",x"B7",x"20",x"4B",x"F7",x"20",x"4C",x"17",x"FF",x"12",x"17",x"FF",x"1B",x"24",x"08",x"8D",
    x"25",x"8D",x"05",x"26",x"F5",x"03",x"78",x"39",x"34",x"04",x"DC",x"90",x"30",x"8B",x"B6",x"20",
    x"4C",x"81",x"10",x"26",x"06",x"7F",x"20",x"4C",x"7C",x"20",x"4B",x"7C",x"20",x"4C",x"B6",x"20",
    x"4B",x"B1",x"22",x"1F",x"35",x"84",x"34",x"06",x"BF",x"20",x"4F",x"B6",x"22",x"19",x"81",x"03",
    x"27",x"04",x"3F",x"26",x"20",x"25",x"F6",x"20",x"4C",x"34",x"04",x"6F",x"E2",x"B6",x"20",x"4B",
    x"C6",x"10",x"3D",x"E3",x"E0",x"58",x"49",x"10",x"83",x"01",x"90",x"23",x"03",x"83",x"01",x"91",
    x"FD",x"20",x"4C",x"BD",x"A0",x"25",x"35",x"04",x"F7",x"20",x"4C",x"10",x"25",x"F5",x"7C",x"35",
    x"86",x"7D",x"22",x"4A",x"27",x"14",x"34",x"04",x"D6",x"F6",x"8D",x"22",x"D6",x"F7",x"8D",x"1E",
    x"D6",x"FD",x"F7",x"22",x"B0",x"7F",x"22",x"4A",x"35",x"04",x"10",x"DE",x"75",x"C1",x"47",x"27",
    x"07",x"C1",x"48",x"27",x"03",x"BD",x"EF",x"81",x"BD",x"EF",x"50",x"7E",x"B0",x"7B",x"2B",x"0F",
    x"BD",x"B4",x"64",x"6F",x"84",x"E6",x"01",x"F7",x"20",x"49",x"BD",x"B3",x"5C",x"6F",x"84",x"39",
    x"BD",x"B2",x"7A",x"25",x"FA",x"30",x"88",x"78",x"CE",x"BD",x"E8",x"C6",x"06",x"A6",x"80",x"A1",
    x"C0",x"26",x"EC",x"5A",x"26",x"F7",x"3F",x"A8",x"42",x"41",x"53",x"49",x"43",x"32",x"88",x"7F",
    x"00",x"00",x"88",x"00",x"00",x"00",x"BD",x"BF",x"49",x"5F",x"20",x"37",x"BD",x"C0",x"48",x"03",
    x"56",x"03",x"62",x"20",x"06",x"8E",x"D1",x"91",x"BD",x"C0",x"48",x"5D",x"10",x"27",x"03",x"E2",
    x"8E",x"21",x"59",x"1F",x"89",x"4D",x"26",x"01",x"39",x"D0",x"4E",x"27",x"D9",x"25",x"0A",x"97",
    x"4E",x"96",x"61",x"97",x"56",x"8E",x"21",x"4E",x"50",x"C1",x"F8",x"2F",x"C9",x"4F",x"64",x"01",
    x"BD",x"BF",x"55",x"D6",x"62",x"2A",x"15",x"63",x"01",x"63",x"02",x"63",x"03",x"0D",x"03",x"27",
    x"08",x"63",x"04",x"63",x"05",x"63",x"06",x"63",x"07",x"43",x"89",x"00",x"97",x"63",x"96",x"03",
    x"27",x"10",x"DC",x"54",x"D9",x"60",x"99",x"5F",x"DD",x"54",x"DC",x"52",x"D9",x"5E",x"99",x"5D",
    x"DD",x"52",x"DC",x"50",x"D9",x"5C",x"99",x"5B",x"DD",x"50",x"96",x"4F",x"99",x"5A",x"97",x"4F",
    x"D6",x"62",x"2A",x"57",x"25",x"02",x"8D",x"7A",x"5F",x"96",x"4F",x"26",x"41",x"DE",x"50",x"DF",
    x"4F",x"96",x"63",x"97",x"51",x"CB",x"08",x"96",x"03",x"27",x"12",x"DE",x"52",x"DF",x"51",x"DE",
    x"54",x"DF",x"53",x"96",x"63",x"97",x"55",x"0F",x"63",x"C1",x"40",x"2D",x"DC",x"0F",x"63",x"C1",
    x"20",x"2D",x"D6",x"4F",x"97",x"4E",x"97",x"56",x"39",x"5C",x"08",x"63",x"96",x"03",x"27",x"08",
    x"09",x"55",x"09",x"54",x"09",x"53",x"09",x"52",x"09",x"51",x"09",x"50",x"09",x"4F",x"2A",x"E9",
    x"96",x"4E",x"34",x"04",x"A0",x"E0",x"97",x"4E",x"23",x"D9",x"8C",x"25",x"08",x"08",x"63",x"86",
    x"00",x"97",x"63",x"20",x"16",x"0C",x"4E",x"27",x"4C",x"06",x"4F",x"06",x"50",x"06",x"51",x"96",
    x"03",x"27",x"08",x"06",x"52",x"06",x"53",x"06",x"54",x"06",x"55",x"24",x"04",x"8D",x"17",x"27",
    x"E4",x"39",x"03",x"56",x"03",x"4F",x"03",x"50",x"03",x"51",x"96",x"03",x"27",x"08",x"03",x"52",
    x"03",x"53",x"03",x"54",x"03",x"55",x"96",x"03",x"27",x"10",x"0C",x"55",x"26",x"16",x"0C",x"54",
    x"26",x"12",x"0C",x"53",x"26",x"0E",x"0C",x"52",x"26",x"0A",x"0C",x"51",x"26",x"06",x"0C",x"50",
    x"26",x"02",x"0C",x"4F",x"39",x"C6",x"06",x"7E",x"B0",x"7B",x"8E",x"21",x"0D",x"A6",x"03",x"97",
    x"63",x"96",x"03",x"27",x"0C",x"A6",x"07",x"97",x"63",x"EE",x"05",x"EF",x"06",x"EE",x"03",x"EF",
    x"04",x"EE",x"01",x"EF",x"02",x"96",x"58",x"A7",x"01",x"CB",x"08",x"2F",x"E0",x"96",x"63",x"C0",
    x"08",x"27",x"16",x"67",x"01",x"66",x"02",x"66",x"03",x"0D",x"03",x"27",x"08",x"66",x"04",x"66",
    x"05",x"66",x"06",x"66",x"07",x"46",x"5C",x"26",x"EA",x"39",x"BD",x"C0",x"48",x"27",x"FA",x"BD",
    x"C0",x"6D",x"34",x"20",x"8E",x"00",x"00",x"9F",x"0E",x"9F",x"0F",x"96",x"03",x"27",x"14",x"9F",
    x"11",x"9F",x"13",x"D6",x"55",x"8D",x"2F",x"D6",x"54",x"8D",x"2B",x"D6",x"53",x"8D",x"27",x"D6",
    x"52",x"8D",x"23",x"D6",x"51",x"8D",x"1F",x"D6",x"63",x"F7",x"22",x"90",x"D6",x"50",x"8D",x"16",
    x"D6",x"63",x"F7",x"22",x"8F",x"D6",x"4F",x"8D",x"11",x"D6",x"63",x"F7",x"22",x"8E",x"BD",x"C1",
    x"6F",x"35",x"20",x"7E",x"BE",x"78",x"10",x"27",x"FF",x"70",x"34",x"04",x"31",x"E4",x"6F",x"E2",
    x"96",x"03",x"27",x"26",x"96",x"60",x"3D",x"ED",x"E2",x"E6",x"A4",x"96",x"5F",x"3D",x"EB",x"E0",
    x"89",x"00",x"34",x"06",x"E6",x"A4",x"96",x"5E",x"3D",x"EB",x"E0",x"89",x"00",x"34",x"06",x"E6",
    x"A4",x"96",x"5D",x"3D",x"EB",x"E0",x"89",x"00",x"34",x"06",x"E6",x"A4",x"96",x"5C",x"3D",x"EB",
    x"E0",x"89",x"00",x"34",x"06",x"E6",x"A4",x"96",x"5B",x"3D",x"EB",x"E0",x"89",x"00",x"34",x"06",
    x"E6",x"A4",x"96",x"5A",x"3D",x"EB",x"E0",x"89",x"00",x"34",x"06",x"96",x"10",x"AB",x"63",x"97",
    x"63",x"0D",x"03",x"27",x"1E",x"96",x"14",x"AB",x"67",x"97",x"63",x"96",x"13",x"A9",x"66",x"97",
    x"14",x"96",x"12",x"A9",x"65",x"97",x"13",x"96",x"11",x"A9",x"64",x"97",x"12",x"96",x"10",x"A9",
    x"63",x"97",x"11",x"96",x"0F",x"A9",x"62",x"97",x"10",x"96",x"0E",x"A9",x"61",x"97",x"0F",x"86",
    x"00",x"A9",x"E4",x"97",x"0E",x"32",x"21",x"39",x"A6",x"01",x"97",x"61",x"1F",x"89",x"8A",x"80",
    x"97",x"5A",x"D8",x"56",x"D7",x"62",x"EE",x"02",x"DF",x"5B",x"96",x"03",x"27",x"08",x"EE",x"04",
    x"DF",x"5D",x"EE",x"06",x"DF",x"5F",x"A6",x"84",x"97",x"59",x"D6",x"4E",x"39",x"4D",x"27",x"18",
    x"9B",x"4E",x"46",x"49",x"28",x"12",x"8B",x"80",x"97",x"4E",x"10",x"27",x"FE",x"28",x"96",x"62",
    x"97",x"56",x"39",x"96",x"56",x"43",x"20",x"02",x"32",x"62",x"10",x"2A",x"FE",x"15",x"7E",x"BF",
    x"25",x"BD",x"C2",x"11",x"27",x"0D",x"8B",x"02",x"25",x"F4",x"0F",x"62",x"BD",x"BE",x"13",x"0C",
    x"4E",x"27",x"EB",x"39",x"C6",x"0B",x"7E",x"B0",x"7B",x"BD",x"C2",x"11",x"8E",x"D1",x"B1",x"0F",
    x"62",x"BD",x"C1",x"84",x"20",x"05",x"8E",x"D0",x"EE",x"8D",x"8D",x"27",x"E7",x"00",x"4E",x"8D",
    x"AC",x"0C",x"4E",x"27",x"C9",x"8E",x"21",x"0E",x"C6",x"03",x"96",x"03",x"27",x"02",x"C6",x"07",
    x"D7",x"02",x"C6",x"01",x"96",x"4F",x"91",x"5A",x"26",x"2A",x"96",x"50",x"91",x"5B",x"26",x"24",
    x"96",x"51",x"91",x"5C",x"26",x"1E",x"96",x"03",x"27",x"18",x"96",x"52",x"91",x"5D",x"26",x"14",
    x"96",x"53",x"91",x"5E",x"26",x"0E",x"96",x"54",x"91",x"5F",x"26",x"08",x"96",x"55",x"91",x"60",
    x"26",x"02",x"1A",x"01",x"1F",x"A8",x"59",x"24",x"0A",x"E7",x"80",x"0A",x"02",x"2B",x"56",x"27",
    x"50",x"C6",x"01",x"1F",x"8A",x"25",x"19",x"4F",x"0D",x"03",x"27",x"08",x"08",x"60",x"09",x"5F",
    x"09",x"5E",x"09",x"5D",x"09",x"5C",x"09",x"5B",x"09",x"5A",x"25",x"D8",x"2B",x"A6",x"20",x"D4",
    x"4F",x"0D",x"03",x"27",x"18",x"96",x"60",x"90",x"55",x"97",x"60",x"96",x"5F",x"92",x"54",x"97",
    x"5F",x"96",x"5E",x"92",x"53",x"97",x"5E",x"96",x"5D",x"92",x"52",x"97",x"5D",x"96",x"5C",x"92",
    x"51",x"97",x"5C",x"96",x"5B",x"92",x"50",x"97",x"5B",x"96",x"5A",x"92",x"4F",x"97",x"5A",x"20",
    x"B6",x"C6",x"40",x"20",x"AE",x"56",x"56",x"56",x"D7",x"63",x"8D",x"03",x"7E",x"BE",x"78",x"9E",
    x"0E",x"9F",x"4F",x"96",x"10",x"97",x"51",x"96",x"03",x"27",x"08",x"9E",x"11",x"9F",x"52",x"9E",
    x"13",x"9F",x"54",x"39",x"D6",x"05",x"C1",x"04",x"27",x"0A",x"25",x"1B",x"EE",x"04",x"DF",x"52",
    x"EE",x"06",x"DF",x"54",x"E6",x"01",x"D7",x"56",x"CA",x"80",x"D7",x"4F",x"0F",x"63",x"E6",x"84",
    x"AE",x"02",x"9F",x"50",x"D7",x"4E",x"39",x"AE",x"84",x"9F",x"50",x"39",x"8E",x"21",x"D7",x"20",
    x"0D",x"8E",x"22",x"A1",x"20",x"08",x"8E",x"22",x"99",x"20",x"03",x"8E",x"22",x"91",x"0D",x"03",
    x"27",x"12",x"20",x"08",x"96",x"05",x"81",x"04",x"27",x"0A",x"25",x"1D",x"DE",x"52",x"EF",x"04",
    x"DE",x"54",x"EF",x"06",x"96",x"4E",x"A7",x"84",x"96",x"56",x"8A",x"7F",x"94",x"4F",x"A7",x"01",
    x"96",x"50",x"A7",x"02",x"96",x"51",x"A7",x"03",x"39",x"96",x"50",x"A7",x"84",x"96",x"51",x"A7",
    x"01",x"39",x"96",x"05",x"81",x"04",x"27",x"0A",x"25",x"10",x"9E",x"5D",x"9F",x"52",x"9E",x"5F",
    x"9F",x"54",x"96",x"61",x"97",x"56",x"9E",x"59",x"9F",x"4E",x"9E",x"5B",x"0F",x"63",x"9F",x"50",
    x"39",x"9E",x"50",x"9F",x"5B",x"96",x"05",x"81",x"04",x"27",x"0A",x"25",x"14",x"9E",x"52",x"9F",
    x"5D",x"9E",x"54",x"9F",x"5F",x"96",x"4F",x"97",x"5A",x"96",x"56",x"97",x"61",x"96",x"4E",x"97",
    x"59",x"39",x"D6",x"4E",x"27",x"08",x"D6",x"56",x"59",x"C6",x"FF",x"25",x"01",x"50",x"39",x"96",
    x"4F",x"80",x"80",x"86",x"00",x"97",x"51",x"D7",x"4E",x"97",x"63",x"97",x"56",x"7E",x"BE",x"74",
    x"8D",x"04",x"1D",x"7E",x"CB",x"03",x"BD",x"CB",x"4C",x"24",x"D7",x"D6",x"50",x"9E",x"50",x"27",
    x"DD",x"20",x"D5",x"8D",x"F1",x"2A",x"D7",x"0F",x"56",x"81",x"02",x"26",x"D1",x"7E",x"CC",x"49",
    x"96",x"61",x"8A",x"7F",x"94",x"5A",x"97",x"5A",x"8E",x"21",x"59",x"E6",x"84",x"27",x"B3",x"E6",
    x"01",x"D8",x"56",x"2B",x"B1",x"D6",x"4E",x"E1",x"84",x"26",x"33",x"E6",x"01",x"CA",x"7F",x"D4",
    x"4F",x"E1",x"01",x"26",x"29",x"D6",x"50",x"E1",x"02",x"26",x"23",x"D6",x"51",x"E0",x"03",x"26",
    x"1D",x"0D",x"03",x"27",x"18",x"D6",x"52",x"E1",x"04",x"26",x"13",x"D6",x"53",x"E1",x"05",x"26",
    x"0D",x"D6",x"54",x"E1",x"06",x"26",x"07",x"D6",x"55",x"E0",x"07",x"26",x"01",x"39",x"56",x"D8",
    x"56",x"7E",x"C2",x"38",x"D6",x"4E",x"27",x"6B",x"C0",x"98",x"96",x"03",x"27",x"02",x"C0",x"20",
    x"96",x"56",x"2A",x"05",x"03",x"58",x"BD",x"BE",x"F4",x"8E",x"21",x"4E",x"C1",x"F8",x"2E",x"06",
    x"BD",x"BF",x"49",x"0F",x"58",x"39",x"0F",x"58",x"96",x"56",x"49",x"06",x"4F",x"7E",x"BF",x"55",
    x"BD",x"CB",x"55",x"25",x"4A",x"BD",x"C2",x"32",x"2A",x"07",x"03",x"56",x"8D",x"03",x"7E",x"CC",
    x"44",x"D6",x"4E",x"BD",x"CB",x"4C",x"25",x"37",x"27",x"06",x"97",x"03",x"C1",x"B8",x"20",x"02",
    x"C1",x"98",x"24",x"2B",x"8D",x"AE",x"D7",x"63",x"96",x"56",x"D7",x"56",x"80",x"80",x"86",x"98",
    x"97",x"4E",x"96",x"51",x"D6",x"03",x"27",x"06",x"86",x"B8",x"97",x"4E",x"96",x"55",x"97",x"00",
    x"7E",x"BE",x"74",x"C6",x"0A",x"CE",x"21",x"4E",x"6F",x"C0",x"5A",x"26",x"FB",x"D7",x"63",x"39",
    x"8D",x"65",x"81",x"4F",x"27",x"0A",x"81",x"42",x"27",x"28",x"81",x"48",x"27",x"10",x"31",x"3F",
    x"8D",x"55",x"24",x"3E",x"81",x"38",x"24",x"3A",x"C6",x"03",x"8D",x"24",x"20",x"F2",x"8D",x"47",
    x"25",x"0A",x"81",x"41",x"25",x"2C",x"81",x"47",x"24",x"28",x"80",x"07",x"C6",x"04",x"8D",x"10",
    x"20",x"EC",x"8D",x"33",x"24",x"1C",x"81",x"31",x"22",x"18",x"C6",x"01",x"8D",x"02",x"20",x"F2",
    x"08",x"51",x"09",x"50",x"10",x"25",x"FB",x"9D",x"5A",x"26",x"F5",x"80",x"30",x"9B",x"51",x"97",
    x"51",x"39",x"34",x"20",x"BD",x"CB",x"A9",x"35",x"A0",x"96",x"05",x"81",x"08",x"4A",x"4A",x"4A",
    x"2F",x"04",x"24",x"02",x"1A",x"02",x"39",x"31",x"21",x"A6",x"A4",x"81",x"20",x"27",x"F8",x"81",
    x"3A",x"24",x"04",x"80",x"30",x"80",x"D0",x"39",x"D6",x"81",x"D0",x"82",x"D7",x"81",x"80",x"30",
    x"34",x"02",x"8D",x"D5",x"2A",x"16",x"8E",x"00",x"0A",x"9F",x"5B",x"BD",x"CC",x"04",x"8D",x"C9",
    x"2A",x"1C",x"4F",x"35",x"04",x"DD",x"5B",x"BD",x"CB",x"E2",x"20",x"55",x"24",x"0D",x"8E",x"C9",
    x"A9",x"BD",x"C2",x"7B",x"2B",x"05",x"BD",x"CB",x"62",x"97",x"03",x"BD",x"C0",x"91",x"BD",x"C2",
    x"11",x"35",x"04",x"BD",x"C2",x"52",x"BD",x"CB",x"8F",x"96",x"03",x"27",x"03",x"BD",x"CB",x"62",
    x"BD",x"CB",x"DD",x"20",x"2C",x"86",x"08",x"97",x"03",x"8C",x"86",x"02",x"97",x"05",x"8D",x"99",
    x"8E",x"00",x"00",x"9F",x"56",x"9F",x"4E",x"9F",x"50",x"9F",x"83",x"9F",x"81",x"25",x"99",x"81",
    x"26",x"10",x"27",x"FF",x"1B",x"81",x"2D",x"26",x"04",x"03",x"57",x"20",x"04",x"81",x"2B",x"26",
    x"05",x"BD",x"C3",x"A7",x"25",x"E7",x"81",x"2E",x"27",x"3C",x"81",x"45",x"27",x"10",x"81",x"25",
    x"27",x"50",x"81",x"23",x"27",x"49",x"81",x"21",x"27",x"46",x"80",x"44",x"26",x"47",x"8D",x"34",
    x"BD",x"C3",x"A7",x"25",x"67",x"81",x"C8",x"27",x"0E",x"81",x"2D",x"27",x"0A",x"81",x"C7",x"27",
    x"08",x"81",x"2B",x"27",x"04",x"20",x"07",x"03",x"84",x"BD",x"C3",x"A7",x"25",x"4E",x"0D",x"84",
    x"27",x"23",x"00",x"83",x"20",x"1F",x"03",x"82",x"27",x"1B",x"BD",x"C3",x"99",x"2A",x"B2",x"BD",
    x"CB",x"8F",x"20",x"AD",x"4D",x"10",x"26",x"06",x"E4",x"43",x"97",x"03",x"7E",x"CB",x"5A",x"4F",
    x"8D",x"F2",x"BD",x"C3",x"A7",x"34",x"20",x"96",x"83",x"90",x"81",x"97",x"83",x"27",x"12",x"2A",
    x"09",x"BD",x"C0",x"A9",x"0C",x"83",x"26",x"F9",x"20",x"07",x"BD",x"C0",x"91",x"0A",x"83",x"26",
    x"F9",x"96",x"57",x"2A",x"03",x"BD",x"CC",x"44",x"0F",x"03",x"35",x"A0",x"D6",x"83",x"C1",x"0A",
    x"24",x"0C",x"58",x"58",x"DB",x"83",x"58",x"80",x"30",x"34",x"04",x"AB",x"E0",x"8C",x"86",x"32",
    x"97",x"83",x"20",x"95",x"34",x"22",x"A6",x"E4",x"46",x"CC",x"01",x"06",x"24",x"04",x"C6",x"04",
    x"86",x"04",x"34",x"04",x"5F",x"08",x"51",x"09",x"50",x"59",x"4A",x"26",x"F8",x"5D",x"26",x"0A",
    x"A6",x"E4",x"4A",x"27",x"05",x"10",x"AC",x"62",x"27",x"0C",x"CB",x"30",x"C1",x"3A",x"25",x"02",
    x"CB",x"07",x"E7",x"A0",x"6F",x"A4",x"35",x"04",x"5A",x"27",x"09",x"A6",x"E4",x"46",x"25",x"D0",
    x"86",x"03",x"20",x"CE",x"35",x"92",x"0F",x"7C",x"30",x"22",x"9F",x"D6",x"BD",x"C3",x"99",x"25",
    x"07",x"97",x"03",x"8D",x"03",x"0F",x"03",x"39",x"C6",x"20",x"96",x"7C",x"85",x"08",x"27",x"02",
    x"C6",x"2B",x"34",x"04",x"BD",x"C2",x"56",x"35",x"02",x"34",x"04",x"2A",x"05",x"BD",x"CC",x"44",
    x"86",x"2D",x"BD",x"C7",x"6C",x"9E",x"D6",x"C6",x"30",x"E7",x"80",x"96",x"7C",x"35",x"04",x"10",
    x"2B",x"02",x"24",x"5D",x"26",x"05",x"6F",x"84",x"30",x"1E",x"39",x"8E",x"00",x"00",x"9F",x"81",
    x"BD",x"C3",x"99",x"10",x"2A",x"00",x"91",x"BD",x"C7",x"2B",x"30",x"22",x"86",x"20",x"D6",x"7C",
    x"C5",x"20",x"27",x"08",x"A1",x"84",x"26",x"04",x"86",x"2A",x"A7",x"84",x"E6",x"84",x"34",x"04",
    x"A7",x"80",x"E6",x"84",x"27",x"14",x"C1",x"45",x"27",x"10",x"C1",x"44",x"27",x"0C",x"C1",x"30",
    x"27",x"EE",x"C1",x"2C",x"27",x"EA",x"C1",x"2E",x"26",x"04",x"86",x"30",x"A7",x"82",x"96",x"7C",
    x"85",x"10",x"27",x"04",x"C6",x"24",x"E7",x"82",x"84",x"04",x"35",x"04",x"26",x"02",x"E7",x"82",
    x"9F",x"50",x"39",x"4A",x"97",x"83",x"D6",x"05",x"CE",x"21",x"4E",x"33",x"C5",x"AE",x"C3",x"34",
    x"10",x"C0",x"02",x"26",x"F8",x"96",x"56",x"D6",x"05",x"34",x"06",x"8D",x"4F",x"35",x"06",x"97",
    x"61",x"CE",x"21",x"59",x"35",x"10",x"AF",x"C1",x"C0",x"02",x"26",x"F8",x"D6",x"83",x"53",x"96",
    x"81",x"34",x"04",x"A1",x"E0",x"25",x"74",x"BD",x"C1",x"F2",x"30",x"23",x"9F",x"D6",x"BD",x"C7",
    x"54",x"1F",x"98",x"BD",x"C8",x"03",x"20",x"1D",x"8D",x"64",x"96",x"83",x"C6",x"02",x"D7",x"81",
    x"C6",x"06",x"0D",x"03",x"27",x"02",x"C6",x"10",x"34",x"04",x"AB",x"E0",x"2B",x"A5",x"34",x"04",
    x"A1",x"E0",x"2E",x"05",x"4C",x"97",x"81",x"86",x"01",x"4A",x"97",x"83",x"BD",x"C6",x"AC",x"C6",
    x"FF",x"5C",x"A6",x"82",x"81",x"30",x"27",x"F9",x"81",x"2E",x"27",x"02",x"30",x"01",x"D7",x"81",
    x"6F",x"84",x"D6",x"83",x"27",x"25",x"86",x"2B",x"5D",x"2A",x"03",x"86",x"2D",x"50",x"A7",x"01",
    x"96",x"03",x"27",x"02",x"86",x"FF",x"8B",x"45",x"A7",x"84",x"86",x"2F",x"4C",x"C0",x"0A",x"24",
    x"FB",x"CB",x"3A",x"ED",x"02",x"6F",x"04",x"30",x"04",x"9F",x"D6",x"30",x"22",x"39",x"4F",x"97",
    x"83",x"D6",x"4E",x"8E",x"C9",x"A8",x"86",x"FA",x"0D",x"03",x"27",x"05",x"8E",x"C9",x"AD",x"86",
    x"F6",x"E1",x"80",x"22",x"0B",x"34",x"02",x"BD",x"BF",x"6A",x"35",x"02",x"9B",x"83",x"20",x"DF",
    x"8E",x"C9",x"BA",x"96",x"03",x"27",x"03",x"8E",x"C9",x"C6",x"BD",x"C2",x"85",x"2F",x"07",x"BD",
    x"C0",x"A9",x"0C",x"83",x"20",x"EA",x"8E",x"C9",x"B6",x"96",x"03",x"27",x"03",x"8E",x"C9",x"BE",
    x"BD",x"C2",x"85",x"2E",x"B8",x"BD",x"C0",x"91",x"0A",x"83",x"20",x"EA",x"BD",x"BE",x"05",x"BD",
    x"C2",x"C4",x"0D",x"03",x"27",x"35",x"8E",x"C9",x"52",x"C6",x"80",x"BD",x"C7",x"50",x"96",x"55",
    x"AB",x"06",x"97",x"55",x"96",x"54",x"A9",x"05",x"97",x"54",x"96",x"53",x"A9",x"04",x"97",x"53",
    x"96",x"52",x"A9",x"03",x"97",x"52",x"8D",x"2A",x"28",x"E4",x"30",x"04",x"8D",x"3A",x"8C",x"C9",
    x"98",x"26",x"D8",x"9E",x"53",x"9F",x"4F",x"96",x"55",x"97",x"51",x"8E",x"C9",x"98",x"C6",x"80",
    x"8D",x"5E",x"4F",x"8D",x"0D",x"28",x"FB",x"8D",x"1F",x"8C",x"C9",x"9E",x"26",x"F2",x"30",x"02",
    x"20",x"2C",x"96",x"51",x"A9",x"02",x"97",x"51",x"96",x"50",x"A9",x"01",x"97",x"50",x"96",x"4F",
    x"A9",x"84",x"97",x"4F",x"5C",x"56",x"59",x"39",x"30",x"03",x"24",x"03",x"C0",x"0B",x"50",x"CB",
    x"2F",x"1F",x"98",x"84",x"7F",x"8D",x"45",x"53",x"C4",x"80",x"39",x"8E",x"C9",x"9E",x"8D",x"20",
    x"86",x"2F",x"97",x"0A",x"DC",x"50",x"0C",x"0A",x"DD",x"50",x"A3",x"84",x"24",x"F8",x"30",x"02",
    x"96",x"0A",x"8D",x"28",x"8C",x"C9",x"A8",x"26",x"E5",x"8D",x"05",x"9E",x"D6",x"6F",x"84",x"39",
    x"0A",x"81",x"26",x"0E",x"86",x"2E",x"8D",x"14",x"9E",x"D6",x"30",x"1F",x"9F",x"45",x"0F",x"82",
    x"20",x"12",x"0A",x"82",x"26",x"10",x"86",x"03",x"97",x"82",x"86",x"2C",x"9F",x"0A",x"9E",x"D6",
    x"A7",x"80",x"9F",x"D6",x"9E",x"0A",x"39",x"9F",x"D6",x"BD",x"C3",x"99",x"10",x"2A",x"00",x"B8",
    x"96",x"7C",x"46",x"10",x"25",x"01",x"55",x"8E",x"06",x"03",x"9F",x"81",x"BD",x"C8",x"19",x"96",
    x"7B",x"80",x"05",x"8D",x"6E",x"8D",x"94",x"96",x"7A",x"26",x"04",x"30",x"1F",x"9F",x"D6",x"4A",
    x"8D",x"61",x"BD",x"C5",x"6A",x"4D",x"27",x"08",x"81",x"2A",x"27",x"04",x"1F",x"98",x"8D",x"BC",
    x"4F",x"8D",x"B9",x"30",x"21",x"30",x"01",x"9F",x"0A",x"96",x"46",x"90",x"0B",x"90",x"7B",x"27",
    x"B5",x"A6",x"84",x"81",x"20",x"27",x"EE",x"81",x"2A",x"27",x"EA",x"4F",x"34",x"02",x"A6",x"80",
    x"81",x"2D",x"27",x"F8",x"81",x"2B",x"27",x"F4",x"81",x"24",x"27",x"F0",x"81",x"30",x"26",x"0F",
    x"A6",x"01",x"BD",x"C3",x"AF",x"24",x"08",x"35",x"02",x"A7",x"82",x"26",x"FA",x"20",x"C6",x"A6",
    x"E0",x"26",x"FC",x"9E",x"0A",x"86",x"25",x"A7",x"82",x"39",x"34",x"02",x"86",x"30",x"BD",x"C7",
    x"6C",x"35",x"02",x"4A",x"2A",x"F4",x"39",x"96",x"83",x"34",x"04",x"AB",x"E0",x"4C",x"97",x"81",
    x"4C",x"80",x"03",x"24",x"FC",x"8B",x"05",x"97",x"82",x"96",x"7C",x"84",x"40",x"26",x"02",x"97",
    x"82",x"39",x"34",x"02",x"BD",x"C7",x"50",x"35",x"02",x"4A",x"2B",x"0B",x"34",x"02",x"86",x"30",
    x"BD",x"C7",x"6C",x"A6",x"E0",x"26",x"EB",x"39",x"96",x"7C",x"46",x"10",x"25",x"00",x"A0",x"8E",
    x"C9",x"CE",x"BD",x"C2",x"85",x"2B",x"05",x"BD",x"C5",x"16",x"20",x"A9",x"C6",x"06",x"96",x"03",
    x"27",x"02",x"C6",x"10",x"96",x"4E",x"97",x"83",x"27",x"07",x"34",x"04",x"BD",x"C6",x"5E",x"35",
    x"04",x"96",x"83",x"2B",x"1C",x"40",x"9B",x"7B",x"34",x"04",x"A0",x"E0",x"8D",x"95",x"8D",x"97",
    x"BD",x"C6",x"AC",x"96",x"83",x"8D",x"B2",x"96",x"83",x"BD",x"C7",x"50",x"9E",x"D6",x"7E",x"C7",
    x"97",x"96",x"7A",x"27",x"01",x"4A",x"9B",x"83",x"2B",x"01",x"4F",x"34",x"06",x"2A",x"0A",x"34",
    x"02",x"BD",x"C0",x"A9",x"35",x"02",x"4C",x"20",x"F4",x"96",x"83",x"A0",x"E0",x"97",x"83",x"AB",
    x"E4",x"35",x"04",x"2B",x"10",x"96",x"7B",x"34",x"04",x"A0",x"E0",x"90",x"83",x"BD",x"C8",x"03",
    x"BD",x"C8",x"07",x"20",x"17",x"96",x"7B",x"BD",x"C8",x"03",x"BD",x"C7",x"54",x"4F",x"34",x"04",
    x"A0",x"E0",x"90",x"83",x"BD",x"C8",x"03",x"8E",x"00",x"00",x"9F",x"81",x"BD",x"C6",x"AC",x"96",
    x"7A",x"26",x"04",x"9E",x"45",x"9F",x"D6",x"9B",x"83",x"7E",x"C7",x"9F",x"BD",x"CB",x"8F",x"C6",
    x"06",x"96",x"03",x"27",x"02",x"C6",x"10",x"96",x"4E",x"34",x"02",x"34",x"04",x"27",x"03",x"BD",
    x"C6",x"5E",x"96",x"7A",x"27",x"01",x"4A",x"9B",x"7B",x"5F",x"34",x"04",x"D6",x"7C",x"C4",x"04",
    x"35",x"04",x"26",x"01",x"53",x"E7",x"A4",x"AB",x"A4",x"A0",x"E4",x"34",x"02",x"2A",x"0A",x"34",
    x"02",x"BD",x"C0",x"A9",x"35",x"02",x"4C",x"20",x"F4",x"A6",x"E4",x"2B",x"01",x"4F",x"40",x"9B",
    x"7B",x"4C",x"AB",x"A4",x"97",x"81",x"0F",x"82",x"BD",x"C6",x"AC",x"35",x"02",x"BD",x"C8",x"29",
    x"9E",x"D6",x"96",x"7A",x"26",x"02",x"30",x"1F",x"35",x"04",x"A6",x"E0",x"27",x"0A",x"96",x"83",
    x"34",x"04",x"AB",x"E0",x"90",x"7B",x"A0",x"A4",x"1F",x"89",x"BD",x"C6",x"36",x"9E",x"D6",x"7E",
    x"C7",x"A2",x"FC",x"72",x"81",x"5B",x"39",x"80",x"00",x"00",x"5A",x"F3",x"10",x"7A",x"40",x"00",
    x"FF",x"F6",x"E7",x"B1",x"8D",x"60",x"00",x"00",x"00",x"E8",x"D4",x"A5",x"10",x"00",x"FF",x"FF",
    x"E8",x"B7",x"89",x"18",x"00",x"00",x"00",x"02",x"54",x"0B",x"E4",x"00",x"FF",x"FF",x"FF",x"C4",
    x"65",x"36",x"00",x"00",x"00",x"00",x"05",x"F5",x"E1",x"00",x"FF",x"FF",x"FF",x"FF",x"67",x"69",
    x"80",x"00",x"00",x"00",x"00",x"0F",x"42",x"40",x"FE",x"79",x"60",x"00",x"27",x"10",x"27",x"10",
    x"03",x"E8",x"00",x"64",x"00",x"0A",x"00",x"01",x"80",x"94",x"74",x"24",x"00",x"91",x"A2",x"15",
    x"02",x"F9",x"00",x"00",x"00",x"00",x"91",x"43",x"4F",x"F8",x"94",x"74",x"23",x"F7",x"B2",x"63",
    x"5F",x"A9",x"31",x"9F",x"FF",x"FC",x"B6",x"0E",x"1B",x"C9",x"BF",x"03",x"FF",x"FD",x"B6",x"0E",
    x"1B",x"C9",x"BF",x"04",x"00",x"00",x"BD",x"CB",x"55",x"24",x"03",x"BD",x"CB",x"EC",x"8E",x"CA",
    x"27",x"7E",x"CB",x"C1",x"96",x"56",x"34",x"02",x"0F",x"56",x"8E",x"C2",x"C4",x"BD",x"CB",x"9C",
    x"9E",x"50",x"86",x"11",x"34",x"12",x"BD",x"C1",x"F2",x"BD",x"C1",x"B1",x"6A",x"E4",x"68",x"62",
    x"69",x"61",x"24",x"F8",x"20",x"0E",x"8D",x"19",x"68",x"62",x"69",x"61",x"24",x"06",x"8E",x"22",
    x"A1",x"BD",x"BF",x"6A",x"6A",x"E4",x"26",x"EE",x"32",x"63",x"A6",x"E0",x"10",x"2B",x"F6",x"96",
    x"39",x"BD",x"C2",x"11",x"7E",x"CB",x"FF",x"10",x"27",x"06",x"2D",x"4D",x"26",x"09",x"96",x"56",
    x"10",x"2B",x"F6",x"70",x"7E",x"BE",x"A4",x"BD",x"C1",x"B1",x"BD",x"C3",x"01",x"8E",x"22",x"A1",
    x"96",x"61",x"BD",x"C2",x"85",x"1F",x"A9",x"26",x"06",x"96",x"4E",x"81",x"90",x"25",x"95",x"6F",
    x"E2",x"96",x"61",x"2A",x"09",x"1F",x"9A",x"26",x"05",x"43",x"D6",x"00",x"E7",x"E4",x"97",x"61",
    x"BD",x"C1",x"F2",x"BD",x"CF",x"9D",x"8E",x"22",x"A1",x"BD",x"BF",x"6A",x"BD",x"D0",x"55",x"66",
    x"E0",x"24",x"06",x"96",x"4E",x"27",x"02",x"03",x"56",x"39",x"9F",x"64",x"BD",x"C1",x"BB",x"8D",
    x"05",x"8D",x"0B",x"8E",x"22",x"91",x"7E",x"BF",x"6A",x"BD",x"CD",x"23",x"9F",x"64",x"BD",x"C1",
    x"B6",x"9E",x"64",x"E6",x"80",x"D7",x"57",x"9F",x"64",x"8D",x"15",x"34",x"14",x"8D",x"E7",x"35",
    x"14",x"3A",x"34",x"14",x"BD",x"BE",x"08",x"8E",x"22",x"99",x"0A",x"57",x"26",x"EF",x"35",x"94",
    x"C6",x"04",x"0D",x"03",x"27",x"01",x"58",x"39",x"BD",x"CB",x"6D",x"BD",x"C2",x"32",x"2B",x"0C",
    x"27",x"2A",x"BE",x"22",x"8B",x"9F",x"4F",x"B6",x"22",x"8D",x"97",x"51",x"BE",x"CA",x"FF",x"9F",
    x"5A",x"B6",x"CB",x"01",x"97",x"5C",x"BD",x"BF",x"72",x"FC",x"22",x"8F",x"C3",x"B0",x"65",x"FD",
    x"22",x"8C",x"F6",x"22",x"8E",x"C9",x"05",x"96",x"0F",x"FD",x"22",x"8A",x"FC",x"22",x"8A",x"97",
    x"63",x"86",x"80",x"DD",x"4E",x"BE",x"22",x"8C",x"9F",x"50",x"0F",x"56",x"7E",x"BE",x"78",x"40",
    x"E6",x"4D",x"4F",x"DD",x"50",x"20",x"35",x"80",x"04",x"27",x"62",x"22",x"4D",x"4C",x"27",x"31",
    x"8D",x"3A",x"27",x"04",x"25",x"2A",x"97",x"03",x"BD",x"BE",x"05",x"0F",x"03",x"8D",x"36",x"27",
    x"02",x"8D",x"50",x"96",x"4E",x"81",x"90",x"10",x"24",x"F3",x"FA",x"96",x"56",x"34",x"02",x"0F",
    x"56",x"BD",x"C2",x"C4",x"A6",x"E0",x"2A",x"04",x"03",x"50",x"03",x"51",x"86",x"02",x"97",x"05",
    x"39",x"96",x"05",x"81",x"03",x"27",x"F9",x"C6",x"0D",x"7E",x"B0",x"7B",x"96",x"05",x"81",x"03",
    x"27",x"F5",x"81",x"04",x"39",x"96",x"05",x"81",x"04",x"39",x"8D",x"F0",x"22",x"FB",x"27",x"02",
    x"8D",x"2D",x"8E",x"00",x"00",x"9F",x"52",x"9F",x"54",x"86",x"08",x"20",x"D1",x"8D",x"DD",x"27",
    x"E8",x"25",x"1C",x"86",x"04",x"97",x"05",x"96",x"4E",x"27",x"DE",x"96",x"52",x"97",x"63",x"8E",
    x"BE",x"CD",x"20",x"18",x"0F",x"03",x"8D",x"C4",x"27",x"04",x"2B",x"03",x"03",x"03",x"39",x"9E",
    x"50",x"9F",x"4F",x"C6",x"90",x"86",x"04",x"97",x"05",x"8E",x"C2",x"3F",x"96",x"03",x"34",x"02",
    x"0F",x"03",x"AD",x"84",x"35",x"02",x"97",x"03",x"39",x"C6",x"98",x"86",x"04",x"97",x"05",x"4F",
    x"97",x"4F",x"97",x"03",x"1A",x"01",x"7E",x"C2",x"47",x"96",x"05",x"81",x"02",x"27",x"1D",x"32",
    x"62",x"96",x"61",x"98",x"56",x"97",x"62",x"96",x"59",x"D6",x"4E",x"6E",x"84",x"8D",x"1D",x"8E",
    x"BD",x"FF",x"8D",x"E5",x"DC",x"5B",x"93",x"50",x"29",x"F3",x"DD",x"50",x"39",x"8E",x"BE",x"0B",
    x"8D",x"D7",x"DC",x"50",x"D3",x"5B",x"28",x"F2",x"8D",x"02",x"20",x"F1",x"9E",x"50",x"34",x"10",
    x"9E",x"5B",x"8D",x"9D",x"BD",x"C2",x"11",x"35",x"10",x"20",x"96",x"8D",x"29",x"8D",x"ED",x"8E",
    x"BF",x"6D",x"8D",x"B5",x"8D",x"48",x"27",x"D2",x"DC",x"50",x"27",x"D0",x"4D",x"26",x"1B",x"96",
    x"5B",x"3D",x"4D",x"26",x"E6",x"34",x"02",x"34",x"04",x"96",x"5C",x"D6",x"51",x"3D",x"E3",x"E1",
    x"25",x"D9",x"2B",x"0E",x"DD",x"50",x"96",x"62",x"20",x"39",x"D6",x"5B",x"26",x"CD",x"D6",x"5C",
    x"20",x"DF",x"10",x"83",x"80",x"00",x"26",x"C3",x"0D",x"62",x"2B",x"9E",x"DD",x"50",x"BD",x"CB",
    x"8F",x"7E",x"CA",x"73",x"BD",x"CB",x"4C",x"24",x"F8",x"8D",x"1A",x"29",x"F1",x"39",x"96",x"50",
    x"98",x"5B",x"97",x"62",x"8D",x"0B",x"DC",x"5B",x"2A",x"06",x"4F",x"5F",x"93",x"5B",x"DD",x"5B",
    x"39",x"96",x"50",x"2A",x"06",x"4F",x"5F",x"93",x"50",x"DD",x"50",x"39",x"DC",x"50",x"10",x"27",
    x"F4",x"32",x"8D",x"DA",x"86",x"10",x"97",x"4F",x"4F",x"5F",x"20",x"0C",x"93",x"50",x"24",x"06",
    x"D3",x"50",x"1C",x"FE",x"20",x"02",x"1A",x"01",x"09",x"5C",x"09",x"5B",x"59",x"49",x"0A",x"4F",
    x"2A",x"EA",x"DD",x"59",x"DC",x"5B",x"20",x"8C",x"96",x"5B",x"34",x"02",x"8D",x"CE",x"DC",x"59",
    x"44",x"56",x"BD",x"CB",x"03",x"E6",x"E0",x"20",x"BA",x"BD",x"CB",x"55",x"24",x"03",x"BD",x"CB",
    x"EC",x"8E",x"C0",x"BB",x"7E",x"CB",x"C1",x"8E",x"C2",x"70",x"BD",x"CB",x"B9",x"DC",x"50",x"93",
    x"5B",x"27",x"07",x"2E",x"03",x"C6",x"FF",x"39",x"C6",x"01",x"39",x"8E",x"CD",x"58",x"D6",x"61",
    x"BD",x"BF",x"6A",x"BD",x"C2",x"11",x"BD",x"C3",x"01",x"0F",x"62",x"96",x"59",x"D6",x"4E",x"7E",
    x"BD",x"FF",x"BD",x"CB",x"84",x"8E",x"CD",x"50",x"BD",x"BE",x"08",x"BD",x"CB",x"84",x"96",x"4E",
    x"81",x"77",x"25",x"D6",x"8D",x"D5",x"8E",x"CD",x"60",x"BD",x"BD",x"FC",x"96",x"56",x"34",x"02",
    x"2A",x"09",x"BD",x"BE",x"05",x"96",x"56",x"2B",x"05",x"03",x"09",x"BD",x"CA",x"73",x"8E",x"CD",
    x"60",x"BD",x"BE",x"08",x"A6",x"E0",x"2A",x"03",x"BD",x"CA",x"73",x"8E",x"CD",x"68",x"8D",x"03",
    x"7E",x"CA",x"7A",x"0D",x"03",x"27",x"03",x"AE",x"02",x"39",x"AE",x"84",x"39",x"BD",x"CB",x"84",
    x"BD",x"C1",x"BB",x"0F",x"09",x"8D",x"B4",x"BD",x"C1",x"B1",x"8E",x"22",x"91",x"BD",x"C1",x"84",
    x"0F",x"56",x"96",x"09",x"8D",x"06",x"8E",x"22",x"A1",x"7E",x"C0",x"B9",x"34",x"02",x"20",x"BB",
    x"81",x"49",x"0F",x"DA",x"A2",x"21",x"68",x"C2",x"7E",x"22",x"F9",x"83",x"6E",x"4E",x"44",x"15",
    x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CD",x"B5",x"CD",x"6C",x"08",x"7D",x"4E",x"8D",
    x"C3",x"4A",x"BF",x"CC",x"F2",x"80",x"B7",x"BC",x"BB",x"86",x"2C",x"A6",x"6B",x"82",x"74",x"79",
    x"AF",x"4E",x"AC",x"D9",x"E2",x"84",x"F1",x"83",x"A6",x"EE",x"8E",x"B8",x"0E",x"86",x"28",x"3C",
    x"1A",x"42",x"8C",x"86",x"5A",x"87",x"99",x"69",x"66",x"73",x"13",x"AA",x"14",x"87",x"23",x"35",
    x"E3",x"3B",x"AD",x"53",x"6F",x"86",x"A5",x"5D",x"E7",x"31",x"2D",x"F2",x"91",x"83",x"49",x"0F",
    x"DA",x"A2",x"21",x"68",x"C2",x"04",x"86",x"1E",x"D7",x"BA",x"87",x"99",x"26",x"64",x"87",x"23",
    x"34",x"58",x"86",x"A5",x"5D",x"E0",x"83",x"49",x"0F",x"DA",x"BD",x"CB",x"4C",x"25",x"1A",x"27",
    x"03",x"BD",x"CB",x"73",x"96",x"56",x"2A",x"06",x"8E",x"CD",x"EC",x"BD",x"BE",x"08",x"96",x"4E",
    x"81",x"90",x"10",x"22",x"01",x"BF",x"BD",x"C2",x"C4",x"9E",x"50",x"39",x"91",x"00",x"00",x"00",
    x"BD",x"CB",x"84",x"96",x"4E",x"10",x"27",x"F0",x"AB",x"4F",x"D6",x"56",x"34",x"06",x"0F",x"56",
    x"96",x"4E",x"81",x"80",x"23",x"07",x"86",x"02",x"A7",x"E4",x"BD",x"C0",x"B6",x"8E",x"CF",x"21",
    x"BD",x"C2",x"85",x"5A",x"26",x"25",x"6C",x"E4",x"BD",x"C1",x"B6",x"8E",x"CF",x"19",x"BD",x"BF",
    x"6A",x"8E",x"D0",x"EE",x"BD",x"BD",x"FC",x"03",x"56",x"BD",x"C1",x"BB",x"BD",x"D0",x"4F",x"8E",
    x"CF",x"19",x"BD",x"BE",x"08",x"8E",x"22",x"91",x"BD",x"C0",x"B9",x"96",x"56",x"34",x"02",x"0F",
    x"56",x"8E",x"CF",x"29",x"BD",x"C2",x"85",x"35",x"02",x"97",x"56",x"5C",x"27",x"45",x"BD",x"C1",
    x"B1",x"BD",x"CA",x"21",x"BD",x"C1",x"B6",x"8E",x"CE",x"AE",x"BD",x"CA",x"89",x"8E",x"22",x"99",
    x"BD",x"BF",x"6A",x"BD",x"C1",x"AC",x"BD",x"D0",x"4F",x"0D",x"03",x"26",x"08",x"8E",x"CE",x"FD",
    x"BD",x"BE",x"08",x"20",x"0C",x"8E",x"CE",x"DC",x"E6",x"80",x"D7",x"57",x"C6",x"08",x"BD",x"CA",
    x"A2",x"8E",x"21",x"D7",x"BD",x"C0",x"B9",x"8E",x"22",x"A1",x"BD",x"BF",x"6A",x"8E",x"22",x"A1",
    x"BD",x"BE",x"08",x"E6",x"E0",x"27",x"10",x"C1",x"01",x"27",x"02",x"03",x"56",x"58",x"58",x"58",
    x"8E",x"CE",x"F9",x"3A",x"BD",x"BE",x"08",x"6D",x"E0",x"2A",x"02",x"03",x"56",x"39",x"CE",x"D3",
    x"CE",x"B2",x"03",x"80",x"D6",x"6B",x"D6",x"CD",x"8C",x"3D",x"E9",x"84",x"87",x"E9",x"FA",x"E4",
    x"6B",x"53",x"1A",x"85",x"A4",x"0B",x"FD",x"CF",x"15",x"E6",x"56",x"84",x"DB",x"05",x"32",x"88",
    x"30",x"E7",x"0E",x"01",x"7C",x"D0",x"86",x"91",x"7F",x"F1",x"10",x"F6",x"04",x"84",x"70",x"62",
    x"4F",x"0A",x"56",x"38",x"83",x"86",x"6E",x"50",x"51",x"90",x"6D",x"1E",x"B4",x"87",x"2C",x"50",
    x"90",x"20",x"5B",x"6D",x"24",x"86",x"24",x"43",x"E5",x"E6",x"24",x"AD",x"4B",x"81",x"34",x"CC",
    x"D3",x"80",x"06",x"0A",x"91",x"C1",x"6B",x"9B",x"2C",x"81",x"49",x"0F",x"DA",x"A2",x"21",x"68",
    x"C2",x"81",x"06",x"0A",x"91",x"C1",x"6B",x"9B",x"2C",x"81",x"5D",x"B3",x"D7",x"42",x"C2",x"65",
    x"53",x"7F",x"09",x"30",x"A2",x"F4",x"F6",x"6A",x"B2",x"65",x"2B",x"CC",x"77",x"11",x"84",x"61",
    x"CF",x"DC",x"50",x"94",x"5B",x"D4",x"5C",x"DD",x"50",x"39",x"DC",x"50",x"9A",x"5B",x"DA",x"5C",
    x"DD",x"50",x"39",x"DC",x"50",x"98",x"5B",x"D8",x"5C",x"DD",x"50",x"39",x"DC",x"50",x"8D",x"F5",
    x"43",x"53",x"DD",x"50",x"39",x"DC",x"50",x"43",x"53",x"8D",x"D8",x"20",x"F3",x"8E",x"CF",x"7B",
    x"BD",x"CB",x"B9",x"DC",x"5B",x"10",x"93",x"50",x"2A",x"02",x"DD",x"50",x"39",x"8E",x"CF",x"7E",
    x"BD",x"CB",x"B9",x"DC",x"5B",x"10",x"93",x"50",x"2A",x"F0",x"39",x"86",x"01",x"8C",x"86",x"FF",
    x"34",x"02",x"BD",x"C2",x"70",x"E1",x"E0",x"26",x"E3",x"8E",x"21",x"59",x"7E",x"C1",x"84",x"8D",
    x"03",x"7E",x"C1",x"BB",x"8E",x"D1",x"91",x"BD",x"BD",x"FC",x"7E",x"CA",x"73",x"BD",x"CB",x"84",
    x"BD",x"C2",x"32",x"2E",x"05",x"C6",x"05",x"7E",x"B0",x"7B",x"96",x"4E",x"80",x"80",x"97",x"D6",
    x"86",x"80",x"97",x"4E",x"8E",x"D1",x"35",x"BD",x"C2",x"85",x"2A",x"06",x"0A",x"D6",x"8D",x"CF",
    x"20",x"0A",x"BD",x"C1",x"B6",x"8D",x"CD",x"8D",x"C6",x"BD",x"D0",x"4F",x"8E",x"D1",x"91",x"8D",
    x"7B",x"BD",x"BE",x"05",x"8E",x"22",x"91",x"BD",x"C0",x"B9",x"8D",x"B5",x"BD",x"CA",x"21",x"0D",
    x"03",x"27",x"0D",x"8E",x"D1",x"03",x"BD",x"CA",x"8C",x"8E",x"22",x"99",x"8D",x"5E",x"20",x"08",
    x"BD",x"C1",x"B6",x"8E",x"D0",x"FA",x"8D",x"54",x"BD",x"C1",x"AC",x"8D",x"52",x"8E",x"D0",x"F6",
    x"BD",x"CD",x"23",x"E6",x"80",x"D7",x"57",x"BD",x"CA",x"B0",x"BD",x"CA",x"A2",x"8E",x"21",x"D7",
    x"BD",x"C0",x"B9",x"8E",x"22",x"91",x"8D",x"34",x"8E",x"22",x"91",x"BD",x"BE",x"08",x"8E",x"D1",
    x"A9",x"8D",x"03",x"8E",x"D1",x"99",x"34",x"10",x"BD",x"C1",x"AC",x"D6",x"D6",x"BD",x"C2",x"52",
    x"BD",x"CA",x"B0",x"1F",x"98",x"BD",x"CB",x"07",x"35",x"10",x"8D",x"10",x"8E",x"21",x"D7",x"7E",
    x"BE",x"08",x"96",x"56",x"2A",x"03",x"7E",x"BE",x"A3",x"7E",x"BF",x"25",x"7E",x"BF",x"6A",x"8E",
    x"22",x"99",x"7E",x"C1",x"84",x"BD",x"CB",x"84",x"BD",x"C1",x"BB",x"8E",x"D0",x"EE",x"0D",x"4E",
    x"27",x"F0",x"8E",x"D1",x"3D",x"8D",x"E5",x"96",x"4E",x"81",x"88",x"24",x"D5",x"BD",x"C3",x"01",
    x"96",x"00",x"4C",x"29",x"CD",x"97",x"D6",x"BD",x"C1",x"B1",x"8E",x"22",x"91",x"8D",x"D3",x"BD",
    x"C3",x"01",x"BD",x"C1",x"B6",x"8E",x"22",x"91",x"BD",x"BD",x"FC",x"8E",x"D1",x"A1",x"CE",x"22",
    x"91",x"8D",x"46",x"8E",x"D1",x"99",x"CE",x"22",x"99",x"8D",x"3E",x"8E",x"22",x"91",x"BD",x"BE",
    x"08",x"BD",x"C1",x"BB",x"BD",x"CA",x"21",x"8E",x"D1",x"49",x"BD",x"CA",x"89",x"BD",x"C1",x"AC",
    x"8D",x"9D",x"8E",x"D1",x"45",x"BD",x"CA",x"89",x"8E",x"22",x"91",x"8D",x"8F",x"8E",x"21",x"D7",
    x"BD",x"C0",x"48",x"BD",x"C1",x"C4",x"BD",x"CB",x"CF",x"8E",x"21",x"D7",x"BD",x"C0",x"B9",x"BD",
    x"BE",x"05",x"96",x"D6",x"9B",x"4E",x"97",x"4E",x"39",x"34",x"50",x"BD",x"C1",x"BB",x"8E",x"22",
    x"A1",x"BD",x"C1",x"84",x"35",x"10",x"BD",x"BF",x"6A",x"35",x"10",x"7E",x"BD",x"FC",x"81",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"D0",x"FE",x"D1",x"1C",x"80",x"8D",x"7E",x"3D",x"01",x"83",
    x"D4",x"3F",x"3A",x"02",x"80",x"CA",x"20",x"AD",x"9A",x"B5",x"E9",x"49",x"85",x"03",x"12",x"51",
    x"00",x"B5",x"7F",x"65",x"87",x"80",x"3F",x"F8",x"95",x"9D",x"AC",x"D2",x"03",x"86",x"8E",x"AC",
    x"02",x"5B",x"3E",x"70",x"78",x"89",x"1C",x"04",x"1F",x"D0",x"A9",x"33",x"EE",x"8A",x"C0",x"5F",
    x"F4",x"E0",x"6C",x"83",x"BC",x"80",x"35",x"04",x"F3",x"33",x"F9",x"DE",x"63",x"81",x"38",x"AA",
    x"3B",x"29",x"5C",x"17",x"F2",x"D1",x"4D",x"D1",x"56",x"D1",x"6F",x"D1",x"78",x"01",x"79",x"08",
    x"53",x"08",x"7F",x"00",x"00",x"00",x"02",x"72",x"04",x"5A",x"21",x"57",x"34",x"90",x"EF",x"79",
    x"78",x"3A",x"5F",x"91",x"50",x"95",x"2B",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",
    x"7C",x"4C",x"BF",x"5B",x"80",x"00",x"00",x"00",x"03",x"6C",x"49",x"9B",x"18",x"67",x"28",x"22",
    x"AA",x"76",x"25",x"78",x"62",x"E1",x"46",x"A6",x"FA",x"7C",x"68",x"B9",x"42",x"8E",x"FE",x"CF",
    x"F5",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"31",x"80",x"00",x"00",x"00",x"00",
    x"00",x"74",x"DE",x"80",x"82",x"E3",x"08",x"65",x"45",x"74",x"DE",x"80",x"82",x"E3",x"08",x"65",
    x"45",x"84",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"BD",x"CB",x"84",x"0D",x"56",x"10",x"2B",
    x"FD",x"E3",x"D6",x"4E",x"26",x"01",x"39",x"4F",x"C5",x"01",x"27",x"08",x"4C",x"5C",x"26",x"04",
    x"C6",x"C0",x"20",x"05",x"C0",x"80",x"57",x"CB",x"80",x"34",x"06",x"C6",x"18",x"0D",x"03",x"27",
    x"02",x"C6",x"38",x"D7",x"02",x"8E",x"21",x"4E",x"CE",x"21",x"0D",x"C6",x"08",x"A6",x"84",x"A7",
    x"0B",x"6F",x"80",x"6F",x"C0",x"5A",x"26",x"F5",x"C6",x"02",x"6D",x"E0",x"26",x"15",x"C6",x"02",
    x"4F",x"0D",x"03",x"27",x"08",x"09",x"60",x"09",x"5F",x"09",x"5E",x"09",x"5D",x"09",x"5C",x"09",
    x"5B",x"09",x"5A",x"0D",x"03",x"27",x"08",x"09",x"14",x"09",x"13",x"09",x"12",x"09",x"11",x"09",
    x"10",x"09",x"0F",x"09",x"0E",x"09",x"0D",x"5A",x"26",x"D6",x"43",x"0D",x"03",x"27",x"08",x"09",
    x"55",x"09",x"54",x"09",x"53",x"09",x"52",x"09",x"51",x"09",x"50",x"09",x"4F",x"09",x"4E",x"9E",
    x"0D",x"9C",x"4E",x"22",x"1C",x"25",x"42",x"9E",x"0F",x"9C",x"50",x"22",x"14",x"25",x"3A",x"0D",
    x"03",x"27",x"0E",x"9E",x"11",x"9C",x"52",x"22",x"08",x"25",x"2E",x"9E",x"13",x"9C",x"54",x"25",
    x"28",x"4F",x"0D",x"03",x"27",x"0E",x"DC",x"13",x"93",x"54",x"DD",x"13",x"DC",x"11",x"D2",x"53",
    x"92",x"52",x"DD",x"11",x"DC",x"0F",x"D2",x"51",x"92",x"50",x"DD",x"0F",x"DC",x"0D",x"D2",x"4F",
    x"92",x"4E",x"DD",x"0D",x"BD",x"BF",x"06",x"20",x"0B",x"8E",x"21",x"51",x"0D",x"03",x"27",x"02",
    x"30",x"04",x"6A",x"84",x"0A",x"02",x"10",x"26",x"FF",x"64",x"04",x"4E",x"06",x"4F",x"06",x"50",
    x"06",x"51",x"06",x"52",x"06",x"53",x"06",x"54",x"06",x"55",x"35",x"02",x"97",x"4E",x"39",x"C6",
    x"02",x"8C",x"C6",x"04",x"8C",x"C6",x"08",x"8D",x"21",x"D7",x"05",x"D1",x"51",x"22",x"5F",x"8E",
    x"23",x"2F",x"7E",x"C1",x"84",x"86",x"02",x"8C",x"86",x"04",x"8C",x"86",x"08",x"BD",x"CB",x"07",
    x"8E",x"23",x"2F",x"BD",x"C1",x"C4",x"D6",x"05",x"20",x"27",x"96",x"05",x"81",x"03",x"27",x"27",
    x"7E",x"CB",x"47",x"8D",x"F5",x"D6",x"51",x"7E",x"CB",x"02",x"8D",x"EE",x"D6",x"51",x"27",x"F7",
    x"10",x"8E",x"23",x"2F",x"4F",x"A7",x"AB",x"7E",x"C4",x"05",x"8D",x"30",x"F7",x"23",x"2F",x"C6",
    x"01",x"D7",x"51",x"86",x"03",x"97",x"05",x"39",x"F6",x"2B",x"69",x"26",x"06",x"3F",x"0A",x"D7",
    x"51",x"27",x"EE",x"7F",x"2B",x"69",x"20",x"E4",x"8D",x"12",x"CB",x"80",x"24",x"DE",x"7E",x"CF",
    x"A5",x"8D",x"09",x"5A",x"C1",x"09",x"22",x"F6",x"CB",x"C0",x"20",x"D0",x"BD",x"CB",x"10",x"DC",
    x"50",x"4D",x"26",x"EA",x"39",x"1F",x"20",x"1F",x"98",x"3F",x"1A",x"C1",x"16",x"26",x"1E",x"3F",
    x"1A",x"4F",x"34",x"06",x"C4",x"F0",x"C1",x"40",x"26",x"04",x"3F",x"1A",x"E7",x"E4",x"35",x"10",
    x"C6",x"99",x"CE",x"D3",x"60",x"AC",x"C1",x"27",x"04",x"5A",x"2B",x"F9",x"5F",x"7E",x"CB",x"02",
    x"41",x"48",x"55",x"48",x"00",x"7B",x"00",x"27",x"00",x"30",x"75",x"48",x"75",x"43",x"75",x"42",
    x"75",x"41",x"6F",x"48",x"6F",x"43",x"6F",x"42",x"6F",x"41",x"69",x"48",x"69",x"43",x"69",x"42",
    x"69",x"41",x"65",x"48",x"65",x"43",x"65",x"42",x"65",x"41",x"61",x"48",x"61",x"43",x"61",x"42",
    x"61",x"41",x"63",x"4B",x"96",x"71",x"27",x"08",x"8E",x"21",x"67",x"BD",x"C1",x"94",x"20",x"0F",
    x"30",x"6E",x"BD",x"C1",x"94",x"E6",x"E8",x"12",x"D7",x"56",x"9E",x"48",x"BD",x"BE",x"08",x"9E",
    x"48",x"BD",x"C1",x"D4",x"30",x"E8",x"13",x"7E",x"C2",x"7B",x"5F",x"34",x"04",x"BD",x"C3",x"33",
    x"35",x"04",x"C1",x"01",x"27",x"1D",x"22",x"02",x"8D",x"19",x"8D",x"20",x"D3",x"50",x"DD",x"50",
    x"CC",x"40",x"98",x"D7",x"4E",x"D6",x"55",x"3D",x"D3",x"4F",x"DD",x"4F",x"86",x"04",x"97",x"05",
    x"7E",x"BE",x"78",x"0F",x"55",x"1F",x"40",x"93",x"1D",x"7E",x"CB",x"03",x"96",x"27",x"90",x"21",
    x"97",x"55",x"DC",x"25",x"93",x"1F",x"2A",x"04",x"0A",x"55",x"8B",x"40",x"39",x"81",x"4F",x"24",
    x"08",x"81",x"32",x"24",x"06",x"81",x"1B",x"25",x"04",x"86",x"2C",x"80",x"17",x"10",x"8E",x"D4",
    x"C0",x"34",x"36",x"4A",x"2B",x"06",x"E6",x"A0",x"2A",x"FC",x"20",x"F7",x"E6",x"A0",x"E7",x"80",
    x"2A",x"FA",x"C4",x"7F",x"E7",x"1F",x"6F",x"84",x"35",x"B6",x"10",x"8E",x"29",x"5B",x"30",x"04",
    x"8D",x"19",x"27",x"62",x"2B",x"24",x"81",x"3A",x"26",x"0D",x"E6",x"84",x"C1",x"8F",x"27",x"F0",
    x"C1",x"8D",x"27",x"EC",x"8C",x"86",x"21",x"8D",x"43",x"20",x"E5",x"BC",x"2C",x"3E",x"26",x"07",
    x"7F",x"2C",x"3E",x"86",x"FF",x"8D",x"35",x"A6",x"80",x"39",x"CE",x"27",x"66",x"81",x"FF",x"26",
    x"04",x"8D",x"E8",x"33",x"45",x"84",x"7F",x"33",x"4A",x"6D",x"C4",x"27",x"D8",x"A0",x"C4",x"2A",
    x"F6",x"AB",x"C4",x"34",x"10",x"8E",x"2B",x"A7",x"34",x"20",x"10",x"AE",x"41",x"8D",x"92",x"35",
    x"20",x"8C",x"8D",x"08",x"A6",x"80",x"26",x"FA",x"35",x"10",x"20",x"A4",x"10",x"8C",x"2A",x"5A",
    x"24",x"04",x"A7",x"A0",x"6F",x"A4",x"39",x"34",x"14",x"5F",x"A6",x"80",x"81",x"61",x"25",x"06",
    x"81",x"7A",x"22",x"02",x"88",x"20",x"A0",x"A0",x"27",x"F0",x"81",x"80",x"27",x"0F",x"31",x"3F",
    x"A6",x"A0",x"2A",x"FC",x"5C",x"AE",x"61",x"E1",x"E4",x"26",x"DF",x"35",x"94",x"32",x"63",x"39",
    x"EE",x"4E",x"65",x"78",x"74",x"20",x"57",x"69",x"74",x"68",x"6F",x"75",x"74",x"20",x"46",x"6F",
    x"F2",x"53",x"79",x"6E",x"74",x"61",x"78",x"20",x"45",x"72",x"72",x"6F",x"F2",x"52",x"65",x"74",
    x"75",x"72",x"6E",x"20",x"57",x"69",x"74",x"68",x"6F",x"75",x"74",x"20",x"47",x"6F",x"73",x"75",
    x"E2",x"4F",x"75",x"74",x"20",x"4F",x"66",x"20",x"44",x"61",x"74",x"E1",x"49",x"6C",x"6C",x"65",
    x"67",x"61",x"6C",x"20",x"46",x"75",x"6E",x"63",x"74",x"69",x"6F",x"6E",x"20",x"43",x"61",x"6C",
    x"EC",x"4F",x"76",x"65",x"72",x"66",x"6C",x"6F",x"F7",x"4F",x"75",x"74",x"20",x"4F",x"66",x"20",
    x"4D",x"65",x"6D",x"6F",x"72",x"F9",x"55",x"6E",x"64",x"65",x"66",x"69",x"6E",x"65",x"64",x"20",
    x"4C",x"69",x"6E",x"65",x"20",x"4E",x"75",x"6D",x"62",x"65",x"F2",x"53",x"75",x"62",x"73",x"63",
    x"72",x"69",x"70",x"74",x"20",x"4F",x"75",x"74",x"20",x"4F",x"66",x"20",x"52",x"61",x"6E",x"67",
    x"E5",x"44",x"75",x"70",x"6C",x"69",x"63",x"61",x"74",x"65",x"20",x"44",x"65",x"66",x"69",x"6E",
    x"69",x"74",x"69",x"6F",x"EE",x"44",x"69",x"76",x"69",x"73",x"69",x"6F",x"6E",x"20",x"42",x"79",
    x"20",x"5A",x"65",x"72",x"EF",x"49",x"6C",x"6C",x"65",x"67",x"61",x"6C",x"20",x"44",x"69",x"72",
    x"65",x"63",x"F4",x"54",x"79",x"70",x"65",x"20",x"4D",x"69",x"73",x"6D",x"61",x"74",x"63",x"E8",
    x"4F",x"75",x"74",x"20",x"4F",x"66",x"20",x"53",x"74",x"72",x"69",x"6E",x"67",x"20",x"53",x"70",
    x"61",x"63",x"E5",x"53",x"74",x"72",x"69",x"6E",x"67",x"20",x"54",x"6F",x"6F",x"20",x"4C",x"6F",
    x"6E",x"E7",x"D3",x"43",x"61",x"6E",x"27",x"74",x"20",x"43",x"6F",x"6E",x"74",x"69",x"6E",x"75",
    x"E5",x"55",x"6E",x"64",x"65",x"66",x"69",x"6E",x"65",x"64",x"20",x"55",x"73",x"65",x"72",x"20",
    x"46",x"75",x"6E",x"63",x"74",x"69",x"6F",x"EE",x"4E",x"6F",x"20",x"52",x"65",x"73",x"75",x"6D",
    x"E5",x"52",x"65",x"73",x"75",x"6D",x"65",x"20",x"57",x"69",x"74",x"68",x"6F",x"75",x"74",x"20",
    x"45",x"72",x"72",x"6F",x"F2",x"55",x"6E",x"64",x"65",x"66",x"69",x"6E",x"65",x"64",x"20",x"45",
    x"72",x"72",x"6F",x"F2",x"4D",x"69",x"73",x"73",x"69",x"6E",x"67",x"20",x"4F",x"70",x"65",x"72",
    x"61",x"6E",x"E4",x"46",x"6F",x"72",x"20",x"57",x"69",x"74",x"68",x"6F",x"75",x"74",x"20",x"4E",
    x"65",x"78",x"F4",x"43",x"61",x"6E",x"27",x"74",x"20",x"45",x"78",x"69",x"F4",x"44",x"6F",x"20",
    x"57",x"69",x"74",x"68",x"6F",x"75",x"74",x"20",x"4C",x"6F",x"6F",x"F0",x"4C",x"6F",x"6F",x"70",
    x"20",x"57",x"69",x"74",x"68",x"6F",x"75",x"74",x"20",x"44",x"EF",x"42",x"61",x"64",x"20",x"46",
    x"69",x"6C",x"65",x"20",x"4E",x"75",x"6D",x"62",x"65",x"F2",x"42",x"61",x"64",x"20",x"46",x"69",
    x"6C",x"65",x"20",x"4D",x"6F",x"64",x"E5",x"46",x"69",x"6C",x"65",x"20",x"41",x"6C",x"72",x"65",
    x"61",x"64",x"79",x"20",x"4F",x"70",x"65",x"EE",x"44",x"65",x"76",x"69",x"63",x"65",x"20",x"49",
    x"2F",x"4F",x"20",x"45",x"72",x"72",x"6F",x"F2",x"49",x"6E",x"70",x"75",x"74",x"20",x"50",x"61",
    x"73",x"74",x"20",x"45",x"6E",x"E4",x"42",x"61",x"64",x"20",x"46",x"69",x"6C",x"65",x"20",x"44",
    x"65",x"73",x"63",x"72",x"69",x"70",x"74",x"6F",x"F2",x"44",x"69",x"72",x"65",x"63",x"74",x"20",
    x"53",x"74",x"61",x"74",x"65",x"6D",x"65",x"6E",x"74",x"20",x"49",x"6E",x"20",x"46",x"69",x"6C",
    x"E5",x"46",x"69",x"6C",x"65",x"20",x"4E",x"6F",x"74",x"20",x"4F",x"70",x"65",x"EE",x"42",x"61",
    x"64",x"20",x"44",x"61",x"74",x"61",x"20",x"49",x"6E",x"20",x"46",x"69",x"6C",x"E5",x"44",x"65",
    x"76",x"69",x"63",x"65",x"20",x"49",x"6E",x"20",x"55",x"73",x"E5",x"44",x"65",x"76",x"69",x"63",
    x"65",x"20",x"55",x"6E",x"61",x"76",x"61",x"69",x"6C",x"61",x"62",x"6C",x"E5",x"50",x"72",x"6F",
    x"74",x"65",x"63",x"74",x"65",x"64",x"20",x"50",x"72",x"6F",x"67",x"72",x"61",x"ED",x"46",x"69",
    x"6C",x"65",x"20",x"4E",x"6F",x"74",x"20",x"46",x"6F",x"75",x"6E",x"E4",x"44",x"69",x"73",x"6B",
    x"20",x"46",x"75",x"6C",x"EC",x"54",x"6F",x"6F",x"20",x"4D",x"61",x"6E",x"79",x"20",x"4F",x"70",
    x"65",x"6E",x"20",x"44",x"69",x"73",x"6B",x"20",x"46",x"69",x"6C",x"65",x"F3",x"44",x"69",x"72",
    x"65",x"63",x"74",x"6F",x"72",x"79",x"20",x"46",x"75",x"6C",x"EC",x"46",x"69",x"6C",x"65",x"20",
    x"41",x"6C",x"72",x"65",x"61",x"64",x"79",x"20",x"45",x"78",x"69",x"73",x"74",x"F3",x"46",x"69",
    x"65",x"6C",x"64",x"20",x"4F",x"76",x"65",x"72",x"66",x"6C",x"6F",x"F7",x"53",x"74",x"72",x"69",
    x"6E",x"67",x"20",x"46",x"69",x"65",x"6C",x"64",x"65",x"E4",x"42",x"61",x"64",x"20",x"52",x"65",
    x"63",x"6F",x"72",x"64",x"20",x"4E",x"75",x"6D",x"62",x"65",x"F2",x"42",x"61",x"64",x"20",x"46",
    x"69",x"6C",x"65",x"20",x"53",x"74",x"72",x"75",x"63",x"74",x"75",x"72",x"E5",x"4E",x"6F",x"20",
    x"44",x"69",x"73",x"EB",x"44",x"69",x"73",x"6B",x"20",x"57",x"72",x"69",x"74",x"65",x"20",x"50",
    x"72",x"6F",x"74",x"65",x"63",x"74",x"65",x"E4",x"4F",x"75",x"74",x"20",x"4F",x"66",x"20",x"46",
    x"69",x"65",x"6C",x"64",x"20",x"42",x"75",x"66",x"66",x"65",x"72",x"F3",x"45",x"6E",x"64",x"20",
    x"4F",x"66",x"20",x"52",x"65",x"63",x"6F",x"72",x"E4",x"56",x"65",x"72",x"69",x"66",x"69",x"63",
    x"61",x"74",x"69",x"6F",x"6E",x"20",x"46",x"61",x"69",x"6C",x"75",x"72",x"E5",x"55",x"6E",x"72",
    x"65",x"61",x"64",x"61",x"62",x"6C",x"65",x"20",x"44",x"69",x"73",x"6B",x"65",x"74",x"74",x"E5",
    x"C4",x"42",x"61",x"64",x"20",x"50",x"69",x"63",x"74",x"75",x"72",x"E5",x"45",x"4E",x"C4",x"46",
    x"4F",x"D2",x"4E",x"45",x"58",x"D4",x"44",x"41",x"54",x"C1",x"44",x"49",x"CD",x"52",x"45",x"41",
    x"C4",x"4C",x"45",x"D4",x"47",x"CF",x"52",x"55",x"CE",x"49",x"C6",x"52",x"45",x"53",x"54",x"4F",
    x"52",x"C5",x"52",x"45",x"54",x"55",x"52",x"CE",x"52",x"45",x"CD",x"A7",x"53",x"54",x"4F",x"D0",
    x"45",x"4C",x"53",x"C5",x"54",x"52",x"4F",x"CE",x"54",x"52",x"4F",x"46",x"C6",x"44",x"45",x"46",
    x"53",x"54",x"D2",x"44",x"45",x"46",x"49",x"4E",x"D4",x"44",x"45",x"46",x"53",x"4E",x"C7",x"44",
    x"45",x"46",x"44",x"42",x"CC",x"4F",x"CE",x"57",x"41",x"49",x"D4",x"45",x"52",x"52",x"4F",x"D2",
    x"52",x"45",x"53",x"55",x"4D",x"C5",x"41",x"55",x"54",x"CF",x"44",x"45",x"4C",x"45",x"54",x"C5",
    x"4C",x"4F",x"43",x"41",x"54",x"C5",x"43",x"4C",x"D3",x"43",x"4F",x"4E",x"53",x"4F",x"4C",x"C5",
    x"50",x"53",x"45",x"D4",x"4D",x"4F",x"54",x"4F",x"D2",x"53",x"4B",x"49",x"50",x"C6",x"45",x"58",
    x"45",x"C3",x"42",x"45",x"45",x"D0",x"43",x"4F",x"4C",x"4F",x"D2",x"4C",x"49",x"4E",x"C5",x"42",
    x"4F",x"D8",x"55",x"4E",x"4D",x"41",x"53",x"CB",x"41",x"54",x"54",x"52",x"C2",x"44",x"45",x"C6",
    x"50",x"4F",x"4B",x"C5",x"50",x"52",x"49",x"4E",x"D4",x"43",x"4F",x"4E",x"D4",x"4C",x"49",x"53",
    x"D4",x"43",x"4C",x"45",x"41",x"D2",x"49",x"4E",x"54",x"45",x"52",x"56",x"41",x"CC",x"4B",x"45",
    x"D9",x"4E",x"45",x"D7",x"53",x"41",x"56",x"C5",x"4C",x"4F",x"41",x"C4",x"4D",x"45",x"52",x"47",
    x"C5",x"4F",x"50",x"45",x"CE",x"43",x"4C",x"4F",x"53",x"C5",x"49",x"4E",x"50",x"45",x"CE",x"50",
    x"45",x"CE",x"50",x"4C",x"41",x"D9",x"54",x"41",x"42",x"A8",x"54",x"CF",x"53",x"55",x"C2",x"46",
    x"CE",x"53",x"50",x"43",x"A8",x"55",x"53",x"49",x"4E",x"C7",x"55",x"53",x"D2",x"45",x"52",x"CC",
    x"45",x"52",x"D2",x"4F",x"46",x"C6",x"54",x"48",x"45",x"CE",x"4E",x"4F",x"D4",x"53",x"54",x"45",
    x"D0",x"AB",x"AD",x"AA",x"AF",x"DE",x"41",x"4E",x"C4",x"4F",x"D2",x"58",x"4F",x"D2",x"45",x"51",
    x"D6",x"49",x"4D",x"D0",x"4D",x"4F",x"C4",x"C0",x"BE",x"BD",x"BC",x"44",x"53",x"4B",x"49",x"4E",
    x"C9",x"44",x"53",x"4B",x"4F",x"A4",x"4B",x"49",x"4C",x"CC",x"4E",x"41",x"4D",x"C5",x"46",x"49",
    x"45",x"4C",x"C4",x"4C",x"53",x"45",x"D4",x"52",x"53",x"45",x"D4",x"50",x"55",x"D4",x"47",x"45",
    x"D4",x"56",x"45",x"52",x"49",x"46",x"D9",x"44",x"45",x"56",x"49",x"43",x"C5",x"44",x"49",x"D2",
    x"46",x"49",x"4C",x"45",x"D3",x"57",x"52",x"49",x"54",x"C5",x"55",x"4E",x"4C",x"4F",x"41",x"C4",
    x"42",x"41",x"43",x"4B",x"55",x"D0",x"43",x"4F",x"50",x"D9",x"43",x"49",x"52",x"43",x"4C",x"C5",
    x"50",x"41",x"49",x"4E",x"D4",x"52",x"45",x"53",x"45",x"D4",x"52",x"45",x"4E",x"55",x"CD",x"53",
    x"57",x"41",x"D0",x"AA",x"57",x"49",x"4E",x"44",x"4F",x"D7",x"50",x"41",x"54",x"54",x"45",x"52",
    x"CE",x"44",x"CF",x"4C",x"4F",x"4F",x"D0",x"45",x"58",x"49",x"D4",x"49",x"4E",x"4D",x"4F",x"55",
    x"53",x"C5",x"4D",x"4F",x"55",x"53",x"C5",x"43",x"48",x"41",x"49",x"CE",x"43",x"4F",x"4D",x"4D",
    x"4F",x"CE",x"53",x"45",x"41",x"52",x"43",x"C8",x"46",x"57",x"C4",x"54",x"55",x"52",x"54",x"4C",
    x"C5",x"53",x"47",x"CE",x"49",x"4E",x"D4",x"41",x"42",x"D3",x"46",x"52",x"C5",x"53",x"51",x"D2",
    x"4C",x"4F",x"C7",x"45",x"58",x"D0",x"43",x"4F",x"D3",x"53",x"49",x"CE",x"54",x"41",x"CE",x"50",
    x"45",x"45",x"CB",x"4C",x"45",x"CE",x"53",x"54",x"52",x"A4",x"56",x"41",x"CC",x"41",x"53",x"C3",
    x"43",x"48",x"52",x"A4",x"45",x"4F",x"C6",x"43",x"49",x"4E",x"D4",x"43",x"53",x"4E",x"C7",x"43",
    x"44",x"42",x"CC",x"46",x"49",x"D8",x"48",x"45",x"58",x"A4",x"4F",x"43",x"54",x"A4",x"53",x"54",
    x"49",x"43",x"CB",x"53",x"54",x"52",x"49",x"C7",x"47",x"52",x"A4",x"4C",x"45",x"46",x"54",x"A4",
    x"52",x"49",x"47",x"48",x"54",x"A4",x"4D",x"49",x"44",x"A4",x"49",x"4E",x"53",x"54",x"D2",x"56",
    x"41",x"52",x"50",x"54",x"D2",x"52",x"4E",x"C4",x"49",x"4E",x"4B",x"45",x"59",x"A4",x"49",x"4E",
    x"50",x"55",x"D4",x"43",x"53",x"52",x"4C",x"49",x"CE",x"50",x"4F",x"49",x"4E",x"D4",x"53",x"43",
    x"52",x"45",x"45",x"CE",x"50",x"4F",x"D3",x"50",x"54",x"52",x"49",x"C7",x"44",x"53",x"4B",x"C6",
    x"43",x"56",x"C9",x"43",x"56",x"D3",x"43",x"56",x"C4",x"4D",x"4B",x"49",x"A4",x"4D",x"4B",x"53",
    x"A4",x"4D",x"4B",x"44",x"A4",x"4C",x"4F",x"C3",x"4C",x"4F",x"C6",x"53",x"50",x"41",x"43",x"45",
    x"A4",x"53",x"54",x"52",x"49",x"4E",x"47",x"A4",x"44",x"53",x"4B",x"49",x"A4",x"46",x"4B",x"45",
    x"59",x"A4",x"4D",x"49",x"4E",x"A8",x"4D",x"41",x"58",x"A8",x"41",x"54",x"CE",x"43",x"52",x"55",
    x"4E",x"43",x"48",x"A4",x"4D",x"54",x"52",x"49",x"C7",x"45",x"56",x"41",x"CC",x"50",x"41",x"4C",
    x"45",x"54",x"54",x"C5",x"42",x"41",x"4E",x"CB",x"48",x"45",x"41",x"C4",x"52",x"4F",x"D4",x"53",
    x"48",x"4F",x"D7",x"5A",x"4F",x"4F",x"CD",x"54",x"52",x"41",x"43",x"C5",x"00",x"34",x"16",x"0D",
    x"DF",x"27",x"1E",x"BD",x"E5",x"4E",x"7D",x"20",x"77",x"2A",x"09",x"F6",x"20",x"1C",x"54",x"25",
    x"03",x"7A",x"A7",x"C0",x"BE",x"20",x"21",x"C6",x"08",x"63",x"84",x"30",x"88",x"D8",x"5A",x"26",
    x"F8",x"35",x"96",x"33",x"3E",x"34",x"70",x"10",x"DF",x"E2",x"86",x"50",x"97",x"9E",x"B6",x"20",
    x"77",x"2B",x"17",x"27",x"13",x"C6",x"7C",x"85",x"01",x"27",x"07",x"C6",x"42",x"BD",x"DD",x"43",
    x"C6",x"50",x"BD",x"DD",x"43",x"BD",x"E3",x"16",x"04",x"9E",x"C6",x"70",x"BD",x"DD",x"43",x"B6",
    x"20",x"1E",x"F6",x"20",x"20",x"DD",x"DA",x"8D",x"42",x"DD",x"D8",x"8D",x"38",x"96",x"DA",x"8D",
    x"34",x"96",x"DB",x"8D",x"30",x"BD",x"DC",x"A6",x"8D",x"93",x"BD",x"DB",x"FE",x"8D",x"8E",x"81",
    x"03",x"27",x"6D",x"81",x"0D",x"27",x"2B",x"BD",x"DD",x"19",x"C6",x"0C",x"8E",x"DE",x"4B",x"EE",
    x"81",x"A1",x"80",x"27",x"0A",x"5A",x"26",x"F7",x"81",x"20",x"25",x"DC",x"CE",x"DC",x"55",x"8D",
    x"0A",x"AD",x"C4",x"20",x"D3",x"4A",x"2B",x"09",x"7E",x"DE",x"37",x"B6",x"20",x"1B",x"F6",x"20",
    x"1C",x"39",x"BD",x"DD",x"C6",x"91",x"D8",x"26",x"02",x"DC",x"D8",x"DD",x"D6",x"BD",x"DD",x"A9",
    x"DD",x"D8",x"DC",x"D6",x"AE",x"E4",x"10",x"93",x"D8",x"22",x"39",x"AC",x"62",x"27",x"35",x"BD",
    x"DE",x"16",x"5D",x"26",x"03",x"BD",x"DD",x"91",x"C1",x"16",x"26",x"0D",x"AC",x"64",x"22",x"24",
    x"E7",x"80",x"DC",x"DD",x"A7",x"80",x"5D",x"27",x"02",x"E7",x"80",x"BD",x"DD",x"D8",x"20",x"D6",
    x"AE",x"E4",x"8D",x"03",x"43",x"35",x"F0",x"6F",x"80",x"BD",x"DC",x"90",x"C6",x"0D",x"8D",x"02",
    x"C6",x"0A",x"3F",x"82",x"8D",x"F1",x"10",x"DE",x"E2",x"7F",x"20",x"2C",x"35",x"F0",x"DE",x"E0",
    x"E6",x"C4",x"27",x"06",x"33",x"41",x"DF",x"E0",x"20",x"07",x"7D",x"22",x"A9",x"26",x"E7",x"3F",
    x"0A",x"D7",x"DC",x"27",x"E9",x"2A",x"1B",x"8E",x"21",x"E4",x"9F",x"E0",x"10",x"8E",x"D8",x"0C",
    x"CE",x"DE",x"ED",x"A6",x"C5",x"2A",x"06",x"10",x"8E",x"D9",x"F1",x"84",x"7F",x"BD",x"D4",x"11",
    x"20",x"CC",x"1F",x"98",x"39",x"FE",x"20",x"5C",x"34",x"40",x"BD",x"DD",x"4B",x"35",x"40",x"FF",
    x"20",x"5C",x"8D",x"2D",x"8D",x"B8",x"C4",x"F0",x"C1",x"40",x"26",x"04",x"8D",x"23",x"8D",x"AE",
    x"BD",x"DB",x"9B",x"20",x"03",x"BD",x"DD",x"4B",x"91",x"D8",x"26",x"06",x"D1",x"D9",x"24",x"02",
    x"D7",x"D9",x"D1",x"9E",x"26",x"0B",x"BD",x"DE",x"45",x"27",x"06",x"8D",x"53",x"91",x"DB",x"27",
    x"04",x"D6",x"DC",x"3F",x"82",x"8D",x"FA",x"BD",x"DE",x"37",x"20",x"34",x"5A",x"26",x"F2",x"91",
    x"DA",x"26",x"EE",x"39",x"8D",x"20",x"8D",x"22",x"D1",x"9E",x"26",x"E5",x"91",x"DB",x"20",x"F1",
    x"BD",x"DD",x"1C",x"BD",x"DD",x"DF",x"8D",x"16",x"C6",x"11",x"8C",x"C6",x"14",x"8C",x"CB",x"40",
    x"20",x"D1",x"03",x"DF",x"26",x"F5",x"0F",x"DF",x"20",x"EE",x"96",x"DA",x"C6",x"01",x"DD",x"D6",
    x"34",x"06",x"C6",x"1F",x"8D",x"BD",x"D6",x"D6",x"8D",x"E4",x"D6",x"D7",x"8D",x"E0",x"35",x"86",
    x"34",x"06",x"B6",x"20",x"59",x"34",x"02",x"BD",x"DD",x"A9",x"91",x"DB",x"22",x"40",x"DD",x"D6",
    x"BD",x"DD",x"C6",x"D6",x"D6",x"91",x"DA",x"25",x"35",x"27",x"12",x"91",x"D8",x"26",x"02",x"0A",
    x"D8",x"6A",x"61",x"33",x"C9",x"FF",x"00",x"8D",x"3B",x"86",x"0A",x"20",x"0B",x"D1",x"DB",x"24",
    x"1D",x"5C",x"D7",x"D6",x"8D",x"2B",x"86",x"0B",x"8D",x"22",x"1F",x"89",x"BD",x"DD",x"9A",x"B6",
    x"20",x"1B",x"4A",x"BD",x"DE",x"40",x"D6",x"DA",x"8D",x"17",x"D6",x"DB",x"8D",x"16",x"EC",x"61",
    x"8D",x"9C",x"35",x"02",x"B7",x"20",x"59",x"35",x"06",x"C6",x"FF",x"21",x"5F",x"F7",x"20",x"2C",
    x"39",x"86",x"20",x"8C",x"86",x"10",x"34",x"02",x"86",x"FF",x"4C",x"C0",x"0A",x"24",x"FB",x"CB",
    x"0A",x"AA",x"E4",x"EA",x"E0",x"34",x"06",x"C6",x"1F",x"8D",x"06",x"35",x"04",x"8D",x"02",x"35",
    x"04",x"3F",x"82",x"34",x"04",x"C6",x"1B",x"8D",x"F8",x"20",x"F4",x"0D",x"DF",x"27",x"D1",x"34",
    x"06",x"8D",x"56",x"91",x"DB",x"26",x"05",x"D1",x"9E",x"26",x"01",x"5A",x"10",x"A3",x"E4",x"10",
    x"25",x"FF",x"5B",x"BD",x"DE",x"45",x"27",x"12",x"1F",x"03",x"5C",x"D1",x"9E",x"26",x"09",x"35",
    x"06",x"BD",x"DC",x"C0",x"DC",x"D6",x"34",x"06",x"1F",x"30",x"10",x"A3",x"E4",x"2B",x"10",x"DD",
    x"D6",x"C6",x"09",x"8D",x"1A",x"DC",x"D6",x"5A",x"26",x"F0",x"D6",x"9E",x"4A",x"20",x"EB",x"32",
    x"62",x"8D",x"04",x"C6",x"20",x"8D",x"AA",x"7E",x"DC",x"B0",x"8D",x"FB",x"7E",x"DC",x"73",x"8D",
    x"F6",x"CE",x"FF",x"FF",x"FF",x"20",x"2E",x"3F",x"82",x"8D",x"34",x"D6",x"9E",x"34",x"06",x"8D",
    x"65",x"C1",x"20",x"35",x"06",x"26",x"20",x"5A",x"26",x"F3",x"4A",x"91",x"DA",x"2D",x"11",x"BD",
    x"DE",x"45",x"26",x"0C",x"20",x"E5",x"BD",x"DB",x"9B",x"4A",x"2B",x"04",x"8D",x"77",x"27",x"F9",
    x"4C",x"5F",x"D1",x"9E",x"27",x"FA",x"5C",x"39",x"DC",x"D6",x"8D",x"F6",x"DD",x"D6",x"39",x"BD",
    x"DB",x"9B",x"4A",x"4C",x"8D",x"5F",x"27",x"FB",x"39",x"C6",x"08",x"D7",x"DC",x"BD",x"DC",x"7C",
    x"BD",x"DB",x"9B",x"34",x"06",x"DD",x"D6",x"8D",x"B0",x"1F",x"01",x"9C",x"D6",x"25",x"36",x"9C",
    x"D6",x"23",x"08",x"8D",x"D3",x"C6",x"08",x"8D",x"96",x"20",x"F4",x"C6",x"20",x"8D",x"8B",x"8D",
    x"26",x"35",x"06",x"7E",x"DC",x"AE",x"34",x"10",x"1F",x"01",x"4F",x"1E",x"01",x"3F",x"1A",x"C1",
    x"16",x"26",x"12",x"0F",x"DE",x"3F",x"1A",x"D7",x"DD",x"C4",x"F0",x"C1",x"40",x"26",x"04",x"3F",
    x"1A",x"D7",x"DE",x"C6",x"16",x"35",x"90",x"8D",x"07",x"63",x"86",x"39",x"91",x"DB",x"27",x"04",
    x"8D",x"03",x"6F",x"86",x"39",x"8E",x"22",x"00",x"6D",x"86",x"39",x"DC",x"7F",x"0B",x"DC",x"8C",
    x"0A",x"DC",x"88",x"09",x"DC",x"7C",x"08",x"DC",x"71",x"18",x"DC",x"35",x"16",x"DC",x"84",x"0C",
    x"DC",x"A2",x"1C",x"DD",x"F3",x"1D",x"DC",x"AA",x"1E",x"DE",x"3C",x"17",x"DD",x"E9",x"7F",x"9D",
    x"2E",x"06",x"A2",x"1D",x"1E",x"2C",x"83",x"99",x"A0",x"28",x"34",x"0B",x"25",x"10",x"22",x"9A",
    x"0A",x"1C",x"2A",x"A4",x"26",x"21",x"03",x"9C",x"05",x"0F",x"1F",x"1B",x"20",x"11",x"24",x"9B",
    x"98",x"08",x"16",x"01",x"2D",x"39",x"8A",x"A1",x"97",x"3B",x"09",x"07",x"9F",x"33",x"2B",x"37",
    x"A6",x"46",x"04",x"3C",x"44",x"32",x"02",x"97",x"02",x"0D",x"02",x"27",x"5C",x"8D",x"08",x"81",
    x"3B",x"27",x"F6",x"8D",x"0F",x"20",x"F2",x"0D",x"02",x"27",x"34",x"A6",x"A0",x"0A",x"02",x"81",
    x"20",x"27",x"F4",x"39",x"81",x"50",x"27",x"62",x"1F",x"89",x"0D",x"02",x"27",x"13",x"8D",x"E7",
    x"8E",x"DF",x"65",x"10",x"A3",x"84",x"27",x"37",x"30",x"03",x"8C",x"DF",x"7A",x"26",x"F4",x"8D",
    x"6B",x"8E",x"DF",x"51",x"E1",x"84",x"27",x"0A",x"30",x"05",x"8C",x"DF",x"65",x"26",x"F5",x"7E",
    x"CF",x"A5",x"8D",x"3D",x"E1",x"01",x"25",x"F7",x"E1",x"02",x"22",x"F3",x"8C",x"DF",x"60",x"26",
    x"05",x"CE",x"DF",x"79",x"E6",x"C5",x"E7",x"98",x"03",x"39",x"8D",x"AB",x"7E",x"C3",x"AF",x"E6",
    x"02",x"0D",x"02",x"27",x"1A",x"8D",x"A0",x"81",x"23",x"26",x"03",x"5C",x"20",x"11",x"81",x"62",
    x"26",x"0B",x"5A",x"C1",x"30",x"22",x"08",x"C6",x"3C",x"8C",x"C6",x"30",x"8C",x"8D",x"1D",x"3F",
    x"9E",x"8D",x"D7",x"24",x"BA",x"5F",x"80",x"30",x"34",x"02",x"86",x"0A",x"3D",x"4D",x"26",x"AF",
    x"EB",x"E0",x"25",x"AB",x"0D",x"02",x"27",x"C1",x"8D",x"C0",x"25",x"EA",x"31",x"3F",x"0C",x"02",
    x"39",x"54",x"01",x"FF",x"20",x"3A",x"41",x"00",x"FF",x"20",x"3D",x"4C",x"01",x"60",x"20",x"3C",
    x"4F",x"01",x"05",x"20",x"3F",x"4F",x"44",x"31",x"45",x"52",x"33",x"49",x"4D",x"35",x"41",x"46",
    x"36",x"4F",x"53",x"38",x"41",x"4C",x"3A",x"49",x"53",x"3C",x"10",x"08",x"04",x"02",x"01",x"8E",
    x"DF",x"8F",x"CE",x"20",x"39",x"C6",x"07",x"A6",x"80",x"A7",x"C0",x"5A",x"26",x"F9",x"39",x"00",
    x"05",x"00",x"18",x"00",x"00",x"02",x"34",x"70",x"8E",x"21",x"D6",x"86",x"19",x"6F",x"80",x"4A",
    x"26",x"FB",x"D6",x"F0",x"1F",x"98",x"3D",x"DD",x"D8",x"0C",x"F1",x"26",x"02",x"0A",x"F1",x"D6",
    x"F1",x"D7",x"DF",x"1F",x"98",x"3D",x"DD",x"E4",x"58",x"49",x"DD",x"DC",x"09",x"DB",x"D6",x"F1",
    x"4F",x"58",x"49",x"83",x"00",x"01",x"34",x"06",x"96",x"D9",x"3D",x"DD",x"E8",x"96",x"D9",x"E6",
    x"E4",x"3D",x"D3",x"E7",x"DD",x"E7",x"96",x"D8",x"E6",x"61",x"3D",x"D3",x"E7",x"DD",x"E7",x"09",
    x"E6",x"96",x"D8",x"E6",x"E1",x"3D",x"D3",x"E6",x"DD",x"E6",x"4F",x"5F",x"93",x"E8",x"DD",x"E8",
    x"DC",x"EA",x"D2",x"E7",x"92",x"E6",x"DD",x"E6",x"4F",x"5F",x"93",x"DE",x"DD",x"DE",x"DC",x"D8",
    x"58",x"49",x"DD",x"D8",x"09",x"D7",x"BD",x"E1",x"C4",x"20",x"03",x"BD",x"E0",x"FF",x"D6",x"DF",
    x"26",x"02",x"35",x"F0",x"96",x"EA",x"2B",x"24",x"0C",x"DF",x"26",x"02",x"0C",x"DE",x"DC",x"EC",
    x"D3",x"E8",x"DD",x"EC",x"DC",x"EA",x"D9",x"E7",x"99",x"E6",x"DD",x"EA",x"DC",x"E8",x"D3",x"D8",
    x"DD",x"E8",x"DC",x"E6",x"D9",x"D7",x"99",x"D6",x"DD",x"E6",x"20",x"CF",x"0D",x"EF",x"27",x"27",
    x"DC",x"A1",x"93",x"DE",x"1F",x"03",x"33",x"5F",x"DC",x"A1",x"D3",x"DE",x"1F",x"01",x"30",x"01",
    x"0D",x"E1",x"27",x"0A",x"DC",x"A3",x"93",x"E0",x"1F",x"02",x"C6",x"FF",x"8D",x"29",x"DC",x"E0",
    x"D3",x"A3",x"1F",x"02",x"5F",x"8D",x"20",x"0C",x"E1",x"DC",x"EC",x"D3",x"E4",x"DD",x"EC",x"DC",
    x"EA",x"D9",x"E3",x"99",x"E2",x"DD",x"EA",x"DC",x"E4",x"D3",x"DC",x"DD",x"E4",x"DC",x"E2",x"D9",
    x"DB",x"99",x"DA",x"DD",x"E2",x"20",x"84",x"0D",x"F2",x"10",x"27",x"05",x"E9",x"96",x"F5",x"91",
    x"F9",x"26",x"10",x"0D",x"EE",x"27",x"07",x"D1",x"F5",x"27",x"08",x"7E",x"E6",x"76",x"D1",x"F5",
    x"27",x"01",x"39",x"34",x"70",x"DC",x"A1",x"40",x"50",x"82",x"00",x"30",x"8B",x"33",x"CB",x"DC",
    x"A3",x"40",x"50",x"82",x"00",x"31",x"AB",x"4F",x"34",x"42",x"1F",x"13",x"BD",x"E1",x"62",x"2B",
    x"18",x"6D",x"E4",x"26",x"11",x"63",x"E4",x"30",x"1F",x"34",x"40",x"AC",x"E1",x"2D",x"02",x"8D",
    x"1C",x"33",x"02",x"30",x"01",x"8C",x"33",x"41",x"8C",x"6F",x"E4",x"30",x"01",x"AC",x"61",x"2F",
    x"DB",x"6D",x"E4",x"2B",x"04",x"30",x"1F",x"8D",x"04",x"32",x"63",x"35",x"F0",x"34",x"70",x"DC",
    x"A1",x"1E",x"13",x"30",x"8B",x"33",x"CB",x"10",x"AE",x"6D",x"BD",x"E6",x"76",x"35",x"F0",x"4F",
    x"5F",x"93",x"E0",x"34",x"06",x"4F",x"5F",x"93",x"DE",x"34",x"06",x"9E",x"DE",x"10",x"9E",x"E0",
    x"8D",x"14",x"9E",x"DE",x"27",x"0E",x"10",x"AE",x"62",x"27",x"09",x"8D",x"09",x"AE",x"E4",x"10",
    x"9E",x"E0",x"8D",x"02",x"35",x"30",x"96",x"F2",x"27",x"04",x"8D",x"36",x"2A",x"51",x"DC",x"A1",
    x"30",x"8B",x"DC",x"A3",x"31",x"AB",x"9C",x"A5",x"25",x"45",x"9C",x"A9",x"22",x"41",x"10",x"9C",
    x"A7",x"25",x"3C",x"10",x"9C",x"AB",x"22",x"37",x"BD",x"E4",x"E9",x"6E",x"9F",x"22",x"84",x"9E",
    x"A1",x"10",x"9E",x"A3",x"7D",x"20",x"36",x"27",x"DD",x"3F",x"90",x"34",x"70",x"8D",x"D7",x"7E",
    x"E4",x"E1",x"34",x"72",x"8E",x"21",x"F3",x"8D",x"0E",x"A7",x"E4",x"8E",x"21",x"F7",x"8D",x"07",
    x"43",x"A4",x"E0",x"98",x"EE",x"35",x"F0",x"A6",x"02",x"A8",x"65",x"2A",x"03",x"A6",x"65",x"39",
    x"EC",x"84",x"EE",x"65",x"8D",x"12",x"EE",x"63",x"34",x"06",x"EC",x"02",x"8D",x"0A",x"A3",x"E1",
    x"26",x"ED",x"6D",x"84",x"2B",x"E7",x"43",x"39",x"34",x"46",x"A8",x"62",x"34",x"01",x"A6",x"61",
    x"2A",x"01",x"50",x"A6",x"64",x"6D",x"63",x"2A",x"01",x"40",x"3D",x"35",x"41",x"2A",x"04",x"40",
    x"50",x"82",x"00",x"35",x"C0",x"8E",x"21",x"F3",x"20",x"03",x"8E",x"21",x"F7",x"86",x"04",x"97",
    x"05",x"7E",x"C1",x"94",x"0D",x"F2",x"27",x"B7",x"8D",x"EB",x"BD",x"CC",x"CB",x"32",x"7C",x"1F",
    x"41",x"BD",x"C1",x"D4",x"8D",x"E4",x"BD",x"CC",x"CB",x"BD",x"C2",x"11",x"1F",x"41",x"BD",x"C1",
    x"94",x"32",x"64",x"BD",x"CC",x"B7",x"5D",x"2B",x"0C",x"03",x"EE",x"8E",x"21",x"F3",x"10",x"8E",
    x"21",x"F7",x"BD",x"E5",x"6F",x"8E",x"21",x"F3",x"8D",x"03",x"8E",x"21",x"F7",x"34",x"10",x"8D",
    x"BC",x"BD",x"CC",x"EB",x"8D",x"12",x"AE",x"E4",x"34",x"40",x"8D",x"B1",x"BD",x"CC",x"E2",x"8D",
    x"07",x"35",x"16",x"EF",x"84",x"ED",x"02",x"39",x"96",x"56",x"34",x"02",x"96",x"4E",x"27",x"04",
    x"8B",x"07",x"97",x"4E",x"BD",x"CB",x"10",x"DE",x"50",x"26",x"07",x"6D",x"E4",x"2A",x"03",x"CE",
    x"FF",x"00",x"35",x"82",x"33",x"84",x"E6",x"C0",x"8D",x"02",x"20",x"FA",x"58",x"8E",x"E2",x"42",
    x"6E",x"95",x"E2",x"83",x"E2",x"7B",x"E2",x"85",x"E2",x"93",x"E2",x"AA",x"E2",x"B0",x"E2",x"B1",
    x"E2",x"B6",x"E2",x"B9",x"E2",x"BE",x"E2",x"C1",x"E2",x"C6",x"E2",x"C9",x"E2",x"CE",x"E2",x"D1",
    x"E2",x"D6",x"E2",x"D9",x"E2",x"E3",x"E2",x"E2",x"E2",x"76",x"E2",x"70",x"E2",x"A5",x"E2",x"9F",
    x"EC",x"C1",x"30",x"CB",x"20",x"07",x"E6",x"C0",x"30",x"C5",x"8C",x"AE",x"C1",x"34",x"40",x"8D",
    x"B3",x"35",x"C0",x"35",x"86",x"A6",x"C0",x"30",x"C4",x"34",x"12",x"8D",x"A7",x"35",x"12",x"4A",
    x"26",x"F7",x"39",x"EC",x"C1",x"34",x"06",x"8D",x"A3",x"35",x"06",x"4A",x"26",x"F7",x"39",x"EC",
    x"C1",x"30",x"CB",x"20",x"07",x"E6",x"C0",x"30",x"C5",x"8C",x"AE",x"C1",x"BF",x"22",x"7D",x"39",
    x"86",x"4F",x"B7",x"22",x"89",x"39",x"8D",x"42",x"8C",x"8D",x"34",x"7E",x"E4",x"E3",x"8D",x"3A",
    x"8C",x"8D",x"2C",x"7E",x"E1",x"5B",x"8D",x"32",x"8C",x"8D",x"24",x"7E",x"E4",x"41",x"8D",x"2A",
    x"8C",x"8D",x"1C",x"4F",x"20",x"07",x"8D",x"22",x"8C",x"8D",x"14",x"86",x"FF",x"97",x"EF",x"7E",
    x"E7",x"56",x"86",x"4F",x"97",x"EF",x"0F",x"F2",x"EC",x"C1",x"DD",x"F0",x"7E",x"DF",x"96",x"E6",
    x"C0",x"1D",x"1F",x"01",x"E6",x"C0",x"1D",x"1F",x"02",x"8C",x"37",x"30",x"7D",x"22",x"89",x"26",
    x"08",x"DC",x"A1",x"30",x"8B",x"DC",x"A3",x"31",x"AB",x"39",x"4F",x"F6",x"20",x"77",x"27",x"05",
    x"4C",x"54",x"24",x"FC",x"48",x"39",x"34",x"56",x"96",x"A0",x"48",x"8E",x"E3",x"B8",x"EE",x"86",
    x"8B",x"08",x"AE",x"86",x"0D",x"9F",x"2A",x"04",x"30",x"1F",x"33",x"5F",x"FF",x"22",x"7F",x"BF",
    x"22",x"81",x"8D",x"D6",x"8E",x"E3",x"41",x"AD",x"96",x"BF",x"22",x"84",x"FD",x"22",x"86",x"35",
    x"D6",x"E3",x"6B",x"E3",x"8F",x"E3",x"8F",x"E3",x"8F",x"E3",x"8F",x"B0",x"7B",x"E3",x"53",x"E3",
    x"53",x"E3",x"B1",x"96",x"9F",x"2A",x"01",x"43",x"84",x"0F",x"34",x"02",x"48",x"48",x"48",x"48",
    x"AA",x"E0",x"97",x"AD",x"8E",x"E3",x"FF",x"CC",x"E4",x"20",x"39",x"C6",x"F0",x"96",x"9F",x"2B",
    x"07",x"53",x"48",x"48",x"48",x"48",x"20",x"01",x"43",x"DD",x"AD",x"8E",x"E3",x"FD",x"B6",x"22",
    x"88",x"27",x"08",x"8E",x"E3",x"FF",x"CC",x"00",x"FF",x"DD",x"AD",x"CC",x"E4",x"15",x"39",x"96",
    x"9F",x"2A",x"01",x"43",x"0F",x"AD",x"0F",x"AE",x"44",x"24",x"02",x"03",x"AE",x"44",x"24",x"02",
    x"03",x"AD",x"8E",x"E4",x"08",x"B6",x"22",x"88",x"27",x"03",x"8E",x"E3",x"FF",x"CC",x"E4",x"15",
    x"39",x"8E",x"E3",x"FF",x"CC",x"E4",x"26",x"39",x"E3",x"C9",x"E3",x"D1",x"E3",x"D7",x"E3",x"DD",
    x"E3",x"E5",x"E3",x"E7",x"E3",x"EB",x"E3",x"E1",x"43",x"A8",x"C4",x"94",x"B0",x"A8",x"C4",x"39",
    x"43",x"94",x"B0",x"AA",x"C4",x"39",x"43",x"94",x"B0",x"A8",x"C4",x"39",x"43",x"43",x"94",x"B0",
    x"43",x"A4",x"C4",x"39",x"43",x"39",x"43",x"AA",x"C4",x"39",x"43",x"A8",x"C4",x"39",x"7A",x"A7",
    x"C0",x"A6",x"C4",x"94",x"AE",x"9A",x"AD",x"A7",x"C4",x"7C",x"A7",x"C0",x"39",x"8D",x"EF",x"96",
    x"AF",x"AD",x"9F",x"22",x"7F",x"A7",x"C4",x"39",x"7A",x"A7",x"C0",x"B6",x"22",x"7C",x"8D",x"F1",
    x"7C",x"A7",x"C0",x"20",x"EA",x"04",x"B0",x"24",x"06",x"86",x"80",x"97",x"B0",x"33",x"41",x"39",
    x"03",x"B0",x"2B",x"08",x"4F",x"39",x"04",x"B0",x"24",x"0F",x"06",x"B0",x"B6",x"A7",x"C0",x"88",
    x"01",x"B7",x"A7",x"C0",x"44",x"24",x"02",x"33",x"41",x"39",x"7D",x"22",x"7C",x"10",x"27",x"00",
    x"A2",x"34",x"70",x"7D",x"20",x"36",x"27",x"0C",x"3F",x"10",x"9E",x"A1",x"10",x"9E",x"A3",x"3F",
    x"0E",x"7E",x"E4",x"E1",x"9F",x"D6",x"10",x"9F",x"D8",x"BD",x"E5",x"A1",x"26",x"F3",x"86",x"28",
    x"97",x"DA",x"DC",x"D8",x"93",x"A3",x"2A",x"06",x"00",x"DA",x"40",x"50",x"82",x"00",x"DD",x"DD",
    x"DC",x"D6",x"93",x"A1",x"2A",x"05",x"BD",x"E5",x"68",x"20",x"E3",x"DD",x"DB",x"9E",x"A1",x"10",
    x"9E",x"A3",x"8D",x"65",x"DC",x"DB",x"10",x"93",x"DD",x"24",x"02",x"DC",x"DD",x"1F",x"02",x"31",
    x"21",x"BE",x"22",x"84",x"44",x"56",x"40",x"50",x"82",x"00",x"DD",x"DF",x"DC",x"DB",x"93",x"DD",
    x"25",x"39",x"DC",x"DD",x"26",x"19",x"BD",x"E6",x"C9",x"20",x"36",x"DC",x"DF",x"D3",x"DD",x"DD",
    x"DF",x"2B",x"08",x"93",x"DB",x"DD",x"DF",x"D6",x"DA",x"33",x"C5",x"AD",x"9F",x"22",x"86",x"AD",
    x"84",x"31",x"3F",x"26",x"E6",x"20",x"1A",x"D6",x"DA",x"33",x"C5",x"DC",x"DF",x"D3",x"DB",x"DD",
    x"DF",x"24",x"08",x"93",x"DD",x"DD",x"DF",x"AD",x"9F",x"22",x"86",x"AD",x"84",x"31",x"3F",x"26",
    x"E6",x"35",x"70",x"9F",x"A1",x"10",x"9F",x"A3",x"39",x"8D",x"48",x"8D",x"2A",x"8D",x"5F",x"1F",
    x"20",x"86",x"28",x"3D",x"1F",x"03",x"B6",x"20",x"77",x"85",x"40",x"27",x"05",x"1F",x"10",x"54",
    x"20",x"0C",x"1F",x"10",x"44",x"56",x"44",x"56",x"54",x"7D",x"20",x"77",x"2A",x"06",x"54",x"24",
    x"03",x"7A",x"A7",x"C0",x"33",x"CB",x"39",x"1F",x"10",x"B6",x"20",x"77",x"85",x"40",x"26",x"0A",
    x"C4",x"07",x"CE",x"E5",x"57",x"A6",x"C5",x"97",x"B0",x"39",x"86",x"F0",x"54",x"24",x"01",x"43",
    x"97",x"B0",x"39",x"86",x"FF",x"F6",x"20",x"77",x"C5",x"40",x"26",x"0D",x"C5",x"01",x"27",x"0B",
    x"34",x"02",x"94",x"AE",x"B7",x"22",x"7C",x"35",x"02",x"94",x"AD",x"97",x"AF",x"39",x"B6",x"A7",
    x"C0",x"8A",x"01",x"B7",x"A7",x"C0",x"39",x"80",x"40",x"20",x"10",x"08",x"04",x"02",x"01",x"FF",
    x"7F",x"3F",x"1F",x"0F",x"07",x"03",x"01",x"00",x"8E",x"21",x"A1",x"10",x"8E",x"21",x"D6",x"34",
    x"46",x"EC",x"84",x"EE",x"A4",x"ED",x"A4",x"EF",x"84",x"EC",x"02",x"EE",x"22",x"ED",x"22",x"EF",
    x"02",x"35",x"C6",x"4F",x"9C",x"A5",x"2C",x"03",x"4C",x"20",x"06",x"9C",x"A9",x"2F",x"02",x"86",
    x"02",x"10",x"9C",x"A7",x"2C",x"03",x"8A",x"04",x"39",x"10",x"9C",x"AB",x"2F",x"02",x"8A",x"08",
    x"39",x"8D",x"E0",x"34",x"02",x"9E",x"A1",x"10",x"9E",x"A3",x"8D",x"D7",x"34",x"02",x"20",x"6E",
    x"A6",x"E4",x"26",x"0A",x"E6",x"61",x"A7",x"61",x"E7",x"E4",x"1F",x"98",x"8D",x"AA",x"84",x"01",
    x"27",x"0F",x"DC",x"A5",x"DD",x"DF",x"DC",x"A1",x"9E",x"D6",x"10",x"9E",x"A3",x"DE",x"D8",x"20",
    x"13",x"A6",x"E4",x"84",x"02",x"27",x"15",x"DC",x"A9",x"DD",x"DF",x"DC",x"D6",x"9E",x"A1",x"10",
    x"9E",x"D8",x"DE",x"A3",x"8D",x"46",x"9F",x"A3",x"DD",x"A1",x"20",x"28",x"A6",x"E4",x"84",x"04",
    x"27",x"0F",x"DC",x"A7",x"DD",x"DF",x"DC",x"A3",x"9E",x"D8",x"10",x"9E",x"A1",x"DE",x"D6",x"20",
    x"0D",x"DC",x"AB",x"DD",x"DF",x"DC",x"D8",x"9E",x"A3",x"10",x"9E",x"D6",x"DE",x"A1",x"8D",x"1C",
    x"9F",x"A1",x"DD",x"A3",x"9E",x"A1",x"10",x"9E",x"A3",x"BD",x"E5",x"83",x"A7",x"E4",x"A6",x"E4",
    x"A4",x"61",x"26",x"06",x"A6",x"E4",x"AA",x"61",x"26",x"86",x"35",x"86",x"34",x"76",x"9C",x"DF",
    x"26",x"06",x"DC",x"DF",x"1F",x"31",x"20",x"2A",x"10",x"93",x"DF",x"26",x"04",x"1F",x"21",x"20",
    x"21",x"EC",x"64",x"E3",x"66",x"47",x"56",x"1F",x"01",x"EC",x"E4",x"E3",x"62",x"47",x"56",x"10",
    x"93",x"DF",x"27",x"0E",x"2C",x"06",x"AF",x"64",x"ED",x"E4",x"20",x"E5",x"AF",x"66",x"ED",x"62",
    x"20",x"DF",x"32",x"68",x"39",x"34",x"40",x"FE",x"22",x"7D",x"1F",x"20",x"C4",x"07",x"53",x"A6",
    x"C5",x"BD",x"E5",x"35",x"35",x"C0",x"B6",x"20",x"36",x"27",x"09",x"3F",x"10",x"1E",x"31",x"3F",
    x"0E",x"1E",x"13",x"39",x"8D",x"DF",x"34",x"70",x"AC",x"64",x"2F",x"02",x"1E",x"13",x"10",x"9C",
    x"A7",x"2D",x"2E",x"10",x"9C",x"AB",x"2E",x"29",x"9C",x"A9",x"2E",x"25",x"9C",x"A5",x"2C",x"02",
    x"9E",x"A5",x"11",x"93",x"A5",x"2D",x"1A",x"11",x"93",x"A9",x"2F",x"02",x"DE",x"A9",x"1F",x"30",
    x"34",x"10",x"A3",x"E1",x"25",x"0B",x"34",x"06",x"BD",x"E4",x"EB",x"35",x"20",x"31",x"21",x"8D",
    x"08",x"35",x"F0",x"AD",x"9F",x"22",x"86",x"25",x"09",x"AD",x"9F",x"22",x"84",x"31",x"3F",x"26",
    x"F2",x"39",x"BE",x"22",x"81",x"B6",x"20",x"77",x"27",x"17",x"2B",x"34",x"85",x"01",x"26",x"52",
    x"85",x"40",x"26",x"6A",x"20",x"E3",x"31",x"38",x"BD",x"E3",x"EE",x"96",x"AF",x"AD",x"84",x"A7",
    x"C0",x"10",x"8C",x"00",x"08",x"24",x"EF",x"31",x"A4",x"26",x"CE",x"39",x"31",x"30",x"96",x"AF",
    x"AD",x"84",x"A7",x"C4",x"7A",x"A7",x"C0",x"96",x"AF",x"AD",x"84",x"A7",x"C0",x"7C",x"A7",x"C0",
    x"10",x"8C",x"00",x"10",x"24",x"E6",x"20",x"DF",x"31",x"38",x"B6",x"22",x"88",x"26",x"0D",x"7A",
    x"A7",x"C0",x"B6",x"22",x"7C",x"AD",x"84",x"A7",x"C4",x"7C",x"A7",x"C0",x"96",x"AF",x"AD",x"84",
    x"A7",x"C0",x"10",x"8C",x"00",x"08",x"24",x"E0",x"20",x"BD",x"31",x"3C",x"96",x"AF",x"AD",x"84",
    x"A7",x"C4",x"7A",x"A7",x"C0",x"96",x"AF",x"AD",x"84",x"A7",x"C0",x"7C",x"A7",x"C0",x"10",x"8C",
    x"00",x"04",x"24",x"E6",x"20",x"A1",x"34",x"70",x"8D",x"38",x"0D",x"EF",x"27",x"2F",x"AE",x"E4",
    x"9C",x"A1",x"2E",x"08",x"27",x"27",x"DE",x"A1",x"9F",x"A1",x"1F",x"31",x"10",x"AE",x"62",x"10",
    x"9C",x"A3",x"2E",x"07",x"DE",x"A3",x"10",x"9F",x"A3",x"1F",x"32",x"33",x"1F",x"9E",x"A1",x"30",
    x"01",x"20",x"03",x"BD",x"E6",x"76",x"31",x"3F",x"10",x"9C",x"A3",x"2E",x"F6",x"35",x"70",x"7E",
    x"E4",x"E3",x"9E",x"A1",x"10",x"9E",x"A3",x"34",x"30",x"AE",x"66",x"8D",x"0B",x"10",x"AE",x"68",
    x"8D",x"06",x"35",x"10",x"8D",x"02",x"35",x"20",x"34",x"30",x"BD",x"E1",x"4F",x"35",x"30",x"7E",
    x"E4",x"41",x"CC",x"00",x"E6",x"BD",x"BB",x"74",x"10",x"DF",x"E1",x"9E",x"6B",x"32",x"89",x"00",
    x"C8",x"9E",x"A1",x"10",x"9E",x"A3",x"BD",x"E5",x"83",x"4D",x"26",x"24",x"3F",x"14",x"D7",x"E3",
    x"DE",x"6E",x"AF",x"56",x"10",x"AF",x"58",x"4F",x"5F",x"ED",x"5A",x"ED",x"5C",x"ED",x"5E",x"33",
    x"C8",x"EC",x"DF",x"DD",x"5C",x"DD",x"DF",x"DC",x"DF",x"83",x"00",x"01",x"DD",x"DF",x"2C",x"04",
    x"10",x"DE",x"E1",x"39",x"DE",x"DD",x"33",x"4A",x"DF",x"DD",x"AE",x"C4",x"2B",x"E9",x"10",x"AE",
    x"42",x"8D",x"5A",x"9F",x"D6",x"AE",x"C4",x"30",x"01",x"8D",x"44",x"25",x"06",x"3F",x"14",x"D1",
    x"E3",x"27",x"F4",x"30",x"1F",x"9F",x"D8",x"9C",x"D6",x"27",x"CC",x"9E",x"D6",x"30",x"01",x"8D",
    x"4D",x"9C",x"D8",x"25",x"F8",x"9E",x"D6",x"30",x"01",x"DE",x"D8",x"BD",x"E6",x"76",x"DE",x"6E",
    x"33",x"56",x"11",x"93",x"DD",x"25",x"11",x"10",x"AC",x"42",x"26",x"F4",x"EC",x"C4",x"10",x"93",
    x"D6",x"2B",x"ED",x"10",x"93",x"D8",x"22",x"E8",x"CC",x"FF",x"FF",x"ED",x"C4",x"20",x"98",x"9C",
    x"A5",x"2D",x"06",x"9C",x"A9",x"2E",x"02",x"4F",x"39",x"43",x"39",x"30",x"1F",x"8D",x"F0",x"25",
    x"06",x"3F",x"14",x"D1",x"E3",x"27",x"F4",x"C6",x"FF",x"D7",x"DA",x"D7",x"DB",x"39",x"34",x"70",
    x"10",x"9F",x"A3",x"10",x"9C",x"A7",x"23",x"08",x"31",x"3F",x"96",x"DB",x"8D",x"14",x"97",x"DB",
    x"10",x"AE",x"62",x"10",x"9C",x"AB",x"24",x"08",x"31",x"21",x"96",x"DA",x"8D",x"04",x"97",x"DA",
    x"35",x"F0",x"34",x"72",x"0F",x"DC",x"3F",x"14",x"D1",x"E3",x"27",x"02",x"0A",x"DC",x"96",x"DC",
    x"A4",x"E4",x"2B",x"13",x"AA",x"E4",x"27",x"0F",x"DE",x"DD",x"AF",x"C4",x"10",x"AF",x"42",x"0C",
    x"E0",x"26",x"02",x"0C",x"DF",x"8D",x"04",x"96",x"DC",x"35",x"F4",x"DC",x"DD",x"83",x"00",x"0A",
    x"34",x"76",x"DE",x"6E",x"33",x"56",x"11",x"A3",x"E4",x"23",x"0F",x"10",x"AC",x"48",x"26",x"F4",
    x"AC",x"44",x"2B",x"F0",x"AC",x"46",x"22",x"EC",x"20",x"35",x"DE",x"6B",x"33",x"C9",x"00",x"E6",
    x"11",x"93",x"DD",x"10",x"24",x"D2",x"94",x"DE",x"DD",x"EC",x"C4",x"ED",x"56",x"EC",x"42",x"ED",
    x"58",x"EC",x"44",x"ED",x"5A",x"EC",x"46",x"ED",x"5C",x"EC",x"48",x"ED",x"5E",x"DC",x"D6",x"ED",
    x"44",x"DC",x"D8",x"ED",x"46",x"9E",x"A3",x"AF",x"48",x"33",x"56",x"DF",x"DD",x"20",x"07",x"DC",
    x"DF",x"83",x"00",x"01",x"DD",x"DF",x"35",x"F6",x"84",x"80",x"C6",x"7F",x"20",x"04",x"84",x"02",
    x"C6",x"FD",x"34",x"02",x"E4",x"2F",x"EA",x"E0",x"E7",x"2F",x"39",x"A8",x"2F",x"84",x"01",x"27",
    x"F9",x"A8",x"2F",x"A7",x"2F",x"20",x"2B",x"33",x"2E",x"5F",x"4D",x"27",x"02",x"E6",x"C4",x"3A",
    x"1F",x"10",x"E7",x"C4",x"39",x"33",x"2C",x"8D",x"F0",x"7E",x"EA",x"A4",x"33",x"2D",x"8D",x"E9",
    x"5F",x"4D",x"27",x"05",x"2B",x"01",x"53",x"E7",x"C4",x"7E",x"EA",x"A4",x"A6",x"2F",x"84",x"01",
    x"27",x"E2",x"34",x"76",x"CE",x"22",x"7F",x"37",x"16",x"34",x"16",x"CC",x"E3",x"D7",x"8E",x"E3",
    x"EB",x"36",x"16",x"7F",x"20",x"36",x"AE",x"A4",x"9F",x"A1",x"EE",x"22",x"DF",x"A3",x"EC",x"24",
    x"30",x"A8",x"10",x"34",x"06",x"EC",x"84",x"26",x"0A",x"35",x"56",x"BF",x"22",x"7F",x"FF",x"22",
    x"81",x"35",x"F6",x"B7",x"22",x"7C",x"26",x"02",x"30",x"01",x"A6",x"80",x"E6",x"61",x"3D",x"58",
    x"49",x"58",x"49",x"58",x"49",x"58",x"49",x"E6",x"80",x"EB",x"E4",x"E7",x"E4",x"34",x"10",x"8D",
    x"1B",x"DC",x"A1",x"30",x"8B",x"D6",x"E3",x"2A",x"02",x"30",x"01",x"DC",x"A3",x"31",x"AB",x"D6",
    x"E4",x"2A",x"02",x"31",x"21",x"BD",x"E4",x"3A",x"35",x"10",x"20",x"B9",x"34",x"06",x"2A",x"01",
    x"50",x"0F",x"E1",x"C1",x"40",x"25",x"05",x"50",x"CB",x"80",x"0A",x"E1",x"8E",x"EB",x"25",x"A6",
    x"85",x"97",x"DB",x"50",x"CB",x"40",x"E6",x"85",x"D7",x"DD",x"A6",x"E4",x"D6",x"DB",x"27",x"03",
    x"D6",x"DD",x"3D",x"D7",x"E4",x"1F",x"89",x"4F",x"6D",x"61",x"2A",x"0B",x"43",x"53",x"03",x"E4",
    x"0C",x"E4",x"26",x"03",x"C3",x"00",x"01",x"1F",x"02",x"A6",x"E4",x"D6",x"DD",x"27",x"03",x"D6",
    x"DB",x"3D",x"D7",x"E3",x"1F",x"89",x"4F",x"0D",x"E1",x"2A",x"0B",x"43",x"53",x"03",x"E3",x"0C",
    x"E3",x"26",x"03",x"C3",x"00",x"01",x"1F",x"01",x"35",x"86",x"1F",x"10",x"4D",x"27",x"08",x"43",
    x"10",x"26",x"E5",x"71",x"50",x"86",x"80",x"33",x"A4",x"AB",x"2E",x"1E",x"89",x"8D",x"8D",x"A6",
    x"48",x"9B",x"E3",x"A7",x"48",x"24",x"02",x"30",x"01",x"EC",x"46",x"30",x"8B",x"AF",x"46",x"A6",
    x"4B",x"9B",x"E4",x"A7",x"4B",x"24",x"02",x"31",x"21",x"EC",x"49",x"31",x"AB",x"10",x"AF",x"49",
    x"31",x"C4",x"EC",x"A4",x"A3",x"26",x"26",x"0D",x"EC",x"22",x"A3",x"29",x"26",x"07",x"EC",x"2C",
    x"A3",x"24",x"26",x"01",x"39",x"BD",x"E9",x"5C",x"A6",x"2F",x"2A",x"19",x"7F",x"20",x"36",x"33",
    x"A4",x"AE",x"C4",x"10",x"AE",x"42",x"9F",x"A1",x"10",x"9F",x"A3",x"AE",x"46",x"10",x"AE",x"49",
    x"BD",x"E4",x"41",x"31",x"C4",x"EC",x"26",x"ED",x"A4",x"EC",x"29",x"ED",x"22",x"EC",x"2C",x"ED",
    x"24",x"7E",x"E9",x"5C",x"A6",x"2F",x"85",x"02",x"27",x"05",x"BD",x"E9",x"5C",x"20",x"E6",x"39",
    x"33",x"A4",x"8E",x"EA",x"BA",x"C6",x"1B",x"7E",x"DF",x"87",x"00",x"A0",x"00",x"64",x"00",x"10",
    x"00",x"A0",x"80",x"00",x"64",x"80",x"00",x"10",x"00",x"00",x"00",x"0F",x"00",x"1E",x"75",x"0F",
    x"4A",x"1E",x"4A",x"00",x"00",x"34",x"70",x"96",x"51",x"97",x"02",x"C6",x"02",x"D7",x"51",x"D6",
    x"02",x"26",x"08",x"E7",x"80",x"E7",x"80",x"D6",x"51",x"35",x"F0",x"BD",x"DE",x"B7",x"81",x"52",
    x"34",x"01",x"27",x"04",x"81",x"4C",x"26",x"14",x"8D",x"25",x"35",x"01",x"27",x"01",x"50",x"34",
    x"04",x"BD",x"DE",x"B7",x"81",x"55",x"27",x"07",x"81",x"44",x"27",x"07",x"7E",x"CF",x"A5",x"6F",
    x"80",x"0C",x"51",x"8D",x"0A",x"E7",x"80",x"27",x"F3",x"35",x"04",x"E7",x"80",x"20",x"C0",x"BD",
    x"DF",x"31",x"0C",x"51",x"39",x"FF",x"FF",x"FF",x"FE",x"FE",x"FD",x"FC",x"FB",x"FA",x"F9",x"F7",
    x"F6",x"F4",x"F2",x"F0",x"EE",x"EC",x"E9",x"E7",x"E4",x"E1",x"DE",x"DB",x"D7",x"D4",x"D0",x"CD",
    x"C9",x"C5",x"C1",x"BD",x"B9",x"B4",x"B0",x"AB",x"A7",x"A2",x"9D",x"98",x"93",x"8E",x"88",x"83",
    x"7E",x"78",x"73",x"6D",x"67",x"62",x"5C",x"56",x"50",x"4A",x"44",x"3E",x"38",x"32",x"2C",x"25",
    x"1F",x"19",x"13",x"0D",x"06",x"00",x"10",x"9F",x"D6",x"9F",x"D8",x"7D",x"22",x"49",x"26",x"47",
    x"0F",x"DB",x"8D",x"43",x"96",x"DE",x"91",x"70",x"22",x"08",x"25",x"09",x"9E",x"DC",x"9C",x"6E",
    x"25",x"03",x"7E",x"BB",x"7B",x"03",x"DB",x"8D",x"2E",x"9E",x"DC",x"96",x"47",x"BD",x"B0",x"7F",
    x"96",x"DE",x"8D",x"0A",x"44",x"56",x"83",x"00",x"01",x"ED",x"9F",x"21",x"45",x"39",x"34",x"12",
    x"8E",x"00",x"00",x"96",x"70",x"A0",x"E0",x"27",x"07",x"30",x"89",x"3F",x"F8",x"4A",x"26",x"F9",
    x"1F",x"10",x"D3",x"6E",x"A3",x"E1",x"39",x"9E",x"45",x"96",x"47",x"30",x"02",x"9F",x"6B",x"97",
    x"6D",x"B6",x"20",x"77",x"84",x"C0",x"97",x"B1",x"BD",x"EC",x"F0",x"9E",x"6B",x"96",x"6D",x"BD",
    x"B0",x"7F",x"0F",x"E5",x"7D",x"22",x"49",x"10",x"26",x"01",x"75",x"96",x"B1",x"8D",x"4C",x"DC",
    x"D8",x"90",x"D6",x"25",x"02",x"D0",x"D7",x"10",x"25",x"E3",x"BA",x"8D",x"73",x"5C",x"58",x"58",
    x"58",x"DD",x"E3",x"8D",x"1C",x"0D",x"B1",x"26",x"05",x"7D",x"22",x"88",x"27",x"07",x"4F",x"5F",
    x"8D",x"5E",x"9F",x"DC",x"39",x"B6",x"20",x"77",x"10",x"26",x"01",x"87",x"03",x"E5",x"7A",x"A7",
    x"C0",x"34",x"66",x"BD",x"ED",x"A5",x"4F",x"E6",x"C4",x"BD",x"EC",x"DC",x"26",x"03",x"8D",x"2F",
    x"8C",x"8D",x"4C",x"0D",x"E1",x"26",x"EF",x"8D",x"D5",x"35",x"E6",x"1E",x"89",x"8D",x"33",x"1E",
    x"89",x"39",x"34",x"06",x"0D",x"E5",x"27",x"15",x"C8",x"80",x"C4",x"F0",x"54",x"A6",x"61",x"85",
    x"08",x"26",x"02",x"CA",x"80",x"84",x"07",x"34",x"04",x"AA",x"E0",x"A7",x"61",x"35",x"86",x"8D",
    x"48",x"4C",x"81",x"FF",x"27",x"08",x"E1",x"C4",x"26",x"04",x"0D",x"E1",x"26",x"F1",x"8D",x"D2",
    x"8D",x"C9",x"0D",x"DB",x"27",x"06",x"BD",x"ED",x"16",x"E7",x"80",x"39",x"30",x"01",x"39",x"8D",
    x"BA",x"31",x"E4",x"8D",x"BD",x"34",x"04",x"8D",x"20",x"4C",x"81",x"FF",x"27",x"0A",x"E6",x"C4",
    x"8D",x"5A",x"27",x"04",x"0D",x"E1",x"26",x"EB",x"8D",x"A1",x"34",x"20",x"E6",x"A2",x"8D",x"D2",
    x"4A",x"26",x"F9",x"10",x"EE",x"E4",x"39",x"A7",x"C4",x"33",x"C8",x"28",x"0A",x"E2",x"26",x"F6",
    x"34",x"22",x"0A",x"E1",x"2A",x"05",x"C6",x"4E",x"7E",x"B0",x"7B",x"96",x"E4",x"97",x"E2",x"8D",
    x"07",x"10",x"9F",x"DF",x"33",x"A4",x"35",x"A2",x"10",x"9E",x"DF",x"0D",x"B1",x"27",x"0B",x"B6",
    x"A7",x"C0",x"88",x"01",x"B7",x"A7",x"C0",x"44",x"24",x"02",x"31",x"21",x"39",x"34",x"02",x"AD",
    x"9F",x"22",x"81",x"8D",x"C2",x"5A",x"35",x"82",x"8D",x"BD",x"5A",x"39",x"34",x"26",x"E6",x"C8",
    x"28",x"96",x"E2",x"4A",x"26",x"06",x"8D",x"D0",x"E6",x"A4",x"8D",x"CF",x"E1",x"61",x"35",x"A6",
    x"96",x"6D",x"97",x"DE",x"DC",x"D6",x"34",x"06",x"BD",x"E5",x"4E",x"6A",x"E4",x"E6",x"61",x"58",
    x"86",x"A0",x"3D",x"0D",x"B1",x"27",x"07",x"64",x"E4",x"24",x"03",x"7A",x"A7",x"C0",x"EB",x"E4",
    x"89",x"00",x"ED",x"E4",x"35",x"C0",x"8C",x"9F",x"F7",x"23",x"17",x"34",x"02",x"8E",x"60",x"00",
    x"0C",x"DE",x"96",x"DE",x"BD",x"B0",x"7F",x"35",x"82",x"8D",x"EB",x"A6",x"80",x"39",x"8D",x"E6",
    x"E6",x"80",x"39",x"34",x"06",x"0D",x"E5",x"27",x"15",x"84",x"78",x"48",x"88",x"80",x"E6",x"E4",
    x"A7",x"E4",x"C4",x"87",x"2B",x"02",x"CA",x"08",x"C4",x"0F",x"EA",x"E4",x"E7",x"E4",x"35",x"86",
    x"8D",x"D7",x"97",x"DA",x"8D",x"D3",x"97",x"E3",x"9B",x"D6",x"81",x"28",x"23",x"08",x"0D",x"B1",
    x"27",x"D0",x"81",x"50",x"22",x"CC",x"8D",x"C1",x"34",x"02",x"9B",x"D7",x"81",x"18",x"35",x"02",
    x"22",x"C0",x"4C",x"48",x"48",x"48",x"97",x"E4",x"10",x"8E",x"EC",x"CD",x"0D",x"B1",x"26",x"13",
    x"8D",x"11",x"7D",x"22",x"88",x"26",x"AB",x"7A",x"A7",x"C0",x"31",x"2B",x"B6",x"20",x"77",x"26",
    x"02",x"03",x"E5",x"34",x"66",x"8D",x"0E",x"8D",x"95",x"27",x"12",x"8D",x"8C",x"8D",x"94",x"AD",
    x"A4",x"26",x"FC",x"20",x"F2",x"DF",x"DF",x"DC",x"E3",x"4C",x"DD",x"E1",x"39",x"BD",x"ED",x"2E",
    x"26",x"02",x"35",x"E6",x"BD",x"ED",x"29",x"BD",x"ED",x"33",x"AD",x"A4",x"26",x"F6",x"20",x"D7",
    x"96",x"47",x"BD",x"B0",x"7F",x"DC",x"6B",x"A3",x"9F",x"21",x"45",x"83",x"00",x"01",x"58",x"49",
    x"1F",x"02",x"39",x"34",x"76",x"96",x"8B",x"B7",x"22",x"91",x"B6",x"20",x"48",x"85",x"0A",x"27",
    x"68",x"96",x"89",x"27",x"0C",x"0F",x"89",x"BD",x"B3",x"5C",x"6D",x"84",x"26",x"03",x"BD",x"EF",
    x"67",x"8D",x"77",x"26",x"05",x"BD",x"EE",x"84",x"27",x"4F",x"BD",x"EE",x"BC",x"FC",x"22",x"AC",
    x"C3",x"00",x"01",x"FD",x"22",x"AC",x"ED",x"05",x"B6",x"20",x"4C",x"4A",x"F6",x"22",x"B1",x"5C",
    x"27",x"03",x"5F",x"44",x"56",x"33",x"CB",x"F6",x"20",x"4C",x"5A",x"B6",x"20",x"48",x"81",x"08",
    x"27",x"10",x"A6",x"A5",x"81",x"FF",x"26",x"03",x"BD",x"EE",x"E3",x"1F",x"31",x"FE",x"20",x"4F",
    x"20",x"09",x"86",x"02",x"A7",x"A5",x"A7",x"07",x"BE",x"20",x"4F",x"F6",x"22",x"B1",x"BD",x"DF",
    x"87",x"B6",x"22",x"91",x"BD",x"B0",x"89",x"35",x"F6",x"8D",x"06",x"3F",x"26",x"25",x"12",x"35",
    x"F6",x"34",x"04",x"F6",x"20",x"48",x"C1",x"08",x"26",x"05",x"DA",x"8D",x"F7",x"20",x"48",x"35",
    x"84",x"B6",x"22",x"91",x"BD",x"B0",x"89",x"7E",x"B3",x"0B",x"B6",x"20",x"49",x"F6",x"20",x"4B",
    x"BE",x"22",x"AE",x"20",x"07",x"10",x"A3",x"03",x"27",x"07",x"30",x"08",x"6D",x"84",x"26",x"F5",
    x"39",x"1C",x"FB",x"39",x"7D",x"22",x"B0",x"27",x"3E",x"BE",x"22",x"AE",x"6D",x"84",x"27",x"37",
    x"A6",x"03",x"2B",x"0F",x"30",x"08",x"6D",x"84",x"26",x"F6",x"8D",x"2C",x"6D",x"07",x"27",x"03",
    x"BD",x"EF",x"81",x"B6",x"20",x"49",x"A7",x"03",x"6F",x"07",x"B6",x"20",x"4B",x"A7",x"04",x"8D",
    x"0B",x"CC",x"FF",x"10",x"A7",x"A0",x"5A",x"26",x"FB",x"1C",x"FB",x"39",x"A6",x"02",x"BD",x"B0",
    x"7F",x"10",x"AE",x"84",x"33",x"A8",x"10",x"39",x"34",x"46",x"FE",x"22",x"AE",x"CC",x"FF",x"FF",
    x"20",x"0B",x"10",x"A3",x"45",x"23",x"04",x"EC",x"45",x"1F",x"31",x"33",x"48",x"6D",x"C4",x"26",
    x"F1",x"35",x"C6",x"34",x"76",x"CC",x"02",x"FF",x"20",x"05",x"34",x"76",x"CC",x"08",x"02",x"34",
    x"04",x"8D",x"44",x"B7",x"20",x"48",x"A6",x"04",x"B7",x"20",x"4B",x"A6",x"03",x"B7",x"20",x"49",
    x"8D",x"BA",x"1F",x"31",x"BD",x"EE",x"51",x"4F",x"4C",x"B7",x"20",x"4C",x"E6",x"A0",x"E1",x"E4",
    x"26",x"12",x"C6",x"01",x"E7",x"3F",x"BF",x"20",x"4F",x"3F",x"26",x"24",x"07",x"C6",x"FF",x"E7",
    x"3F",x"7E",x"EE",x"61",x"F6",x"22",x"B1",x"3A",x"5C",x"26",x"02",x"30",x"01",x"81",x"10",x"26",
    x"D7",x"8D",x"0E",x"32",x"61",x"35",x"F6",x"34",x"56",x"8E",x"20",x"48",x"CE",x"22",x"92",x"20",
    x"08",x"34",x"56",x"CE",x"20",x"48",x"8E",x"22",x"92",x"C6",x"09",x"BD",x"DF",x"87",x"35",x"D6",
    x"34",x"16",x"4F",x"5F",x"FD",x"22",x"AC",x"53",x"BE",x"22",x"AE",x"20",x"04",x"E7",x"03",x"30",
    x"08",x"6D",x"84",x"26",x"F8",x"35",x"96",x"34",x"16",x"B6",x"20",x"49",x"C6",x"FF",x"BE",x"22",
    x"AE",x"20",x"08",x"A1",x"03",x"26",x"02",x"E7",x"03",x"30",x"08",x"6D",x"84",x"26",x"F4",x"35",
    x"96",x"34",x"12",x"96",x"8B",x"34",x"02",x"BE",x"22",x"AE",x"20",x"0B",x"6D",x"03",x"2B",x"05",
    x"BD",x"EE",x"EA",x"6F",x"07",x"30",x"08",x"6D",x"84",x"26",x"F1",x"35",x"02",x"BD",x"B0",x"89",
    x"35",x"92",x"34",x"06",x"86",x"10",x"F6",x"22",x"B1",x"5C",x"27",x"01",x"44",x"5F",x"C3",x"00",
    x"10",x"1F",x"03",x"35",x"86",x"B6",x"22",x"19",x"81",x"03",x"26",x"03",x"7F",x"22",x"B0",x"39",
    x"31",x"38",x"2E",x"30",x"39",x"2E",x"38",x"36",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7E",x"B0",x"21",x"B0",x"1A");

  CONSTANT ROM_BASIC6_3 : arr8 := (
    x"1B",x"38",x"34",x"02",x"B6",x"A7",x"C0",x"84",x"DF",x"B7",x"A7",x"C0",x"35",x"02",x"AD",x"C4",
    x"34",x"02",x"B6",x"A7",x"C0",x"8A",x"20",x"B7",x"A7",x"C0",x"A6",x"E0",x"39",x"CE",x"B0",x"26",
    x"20",x"E0",x"CE",x"CB",x"10",x"20",x"DB",x"CE",x"CB",x"07",x"20",x"D6",x"9E",x"48",x"96",x"4A",
    x"BD",x"DC",x"27",x"CE",x"C1",x"C4",x"20",x"CA",x"CE",x"D3",x"08",x"20",x"C5",x"92",x"50",x"93",
    x"01",x"92",x"63",x"12",x"18",x"A1",x"B9",x"9F",x"9D",x"A0",x"55",x"9C",x"E2",x"9C",x"EB",x"9D",
    x"2D",x"51",x"6F",x"A2",x"E3",x"0F",x"89",x"A2",x"EA",x"0E",x"FF",x"A2",x"FA",x"27",x"1C",x"9B",
    x"10",x"9B",x"6D",x"9B",x"5A",x"92",x"F0",x"0F",x"6F",x"0F",x"70",x"29",x"B2",x"29",x"C3",x"A3",
    x"18",x"4E",x"9D",x"4E",x"B9",x"4E",x"A2",x"53",x"91",x"59",x"12",x"4D",x"DE",x"40",x"38",x"67",
    x"4C",x"69",x"AD",x"72",x"1A",x"72",x"21",x"67",x"83",x"69",x"E2",x"38",x"0D",x"A2",x"AF",x"A2",
    x"B2",x"A2",x"B5",x"A2",x"C5",x"A2",x"C8",x"A2",x"CB",x"3A",x"1B",x"3B",x"F4",x"10",x"A3",x"50",
    x"8D",x"77",x"B6",x"A3",x"21",x"4D",x"F7",x"4D",x"F2",x"9D",x"F0",x"11",x"04",x"29",x"CB",x"11",
    x"2C",x"28",x"A2",x"52",x"01",x"7E",x"18",x"7E",x"1E",x"7E",x"2B",x"7E",x"24",x"7E",x"36",x"79",
    x"CB",x"DD",x"79",x"CB",x"CF",x"7C",x"CB",x"FF",x"7C",x"CC",x"A9",x"7F",x"C9",x"D6",x"50",x"CF",
    x"31",x"46",x"CF",x"3A",x"3C",x"CF",x"43",x"32",x"CF",x"4C",x"28",x"CF",x"55",x"7A",x"CC",x"98",
    x"7B",x"CC",x"6C",x"CC",x"B7",x"B5",x"0F",x"E5",x"02",x"E5",x"95",x"B6",x"E4",x"BC",x"B6",x"CE",
    x"0A",x"B7",x"CF",x"B6",x"68",x"B6",x"54",x"B7",x"18",x"B4",x"F4",x"B6",x"B9",x"B6",x"E7",x"B6",
    x"E7",x"B5",x"19",x"B6",x"E7",x"C5",x"F9",x"C6",x"28",x"C5",x"55",x"C5",x"58",x"C5",x"5B",x"C5",
    x"5E",x"DA",x"62",x"C1",x"C1",x"C8",x"C0",x"C8",x"CB",x"C6",x"2F",x"C5",x"99",x"E0",x"B8",x"D9",
    x"A9",x"E1",x"28",x"E2",x"80",x"E0",x"34",x"DF",x"90",x"C2",x"06",x"D9",x"A6",x"E1",x"9C",x"E2",
    x"8A",x"E3",x"77",x"B8",x"F4",x"E0",x"FA",x"C9",x"29",x"C1",x"9F",x"C2",x"6B",x"B5",x"41",x"D1",
    x"9E",x"B5",x"57",x"C9",x"90",x"B8",x"F4",x"B4",x"2C",x"D1",x"DD",x"D4",x"A0",x"D4",x"98",x"D3",
    x"D1",x"D3",x"8B",x"DA",x"A2",x"D9",x"E6",x"E4",x"8F",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",
    x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",
    x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",
    x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",x"F4",x"B8",
    x"F4",x"E9",x"CC",x"E7",x"6C",x"E9",x"C1",x"E9",x"EE",x"EA",x"62",x"C0",x"B8",x"C0",x"B7",x"EB",
    x"D0",x"EB",x"D1",x"E7",x"EA",x"E7",x"FA",x"E8",x"23",x"E9",x"51",x"C3",x"59",x"EC",x"BA",x"EC",
    x"9B",x"EC",x"00",x"E3",x"2E",x"E3",x"F8",x"B1",x"DF",x"CA",x"30",x"BD",x"8C",x"EB",x"CF",x"E3",
    x"80",x"E3",x"CF",x"E6",x"26",x"E6",x"55",x"E6",x"D9",x"DA",x"9A",x"B8",x"F4",x"D7",x"AC",x"D8",
    x"49",x"CC",x"A6",x"EE",x"3F",x"EE",x"C0",x"0D",x"0A",x"42",x"72",x"65",x"61",x"6B",x"00",x"3F",
    x"80",x"4F",x"58",x"D3",x"1D",x"C3",x"00",x"3A",x"25",x"12",x"10",x"DF",x"15",x"93",x"15",x"22",
    x"0B",x"39",x"86",x"11",x"97",x"77",x"BD",x"D3",x"4F",x"0F",x"77",x"39",x"C6",x"07",x"9E",x"28",
    x"30",x"1F",x"9F",x"75",x"8C",x"C6",x"38",x"F7",x"2C",x"26",x"BD",x"27",x"CD",x"BD",x"27",x"D0",
    x"8D",x"E0",x"7F",x"2C",x"45",x"0F",x"03",x"8E",x"00",x"00",x"BF",x"23",x"20",x"9F",x"2A",x"BD",
    x"DF",x"E1",x"DE",x"31",x"FF",x"2C",x"2A",x"30",x"41",x"27",x"03",x"FF",x"2C",x"40",x"B6",x"29",
    x"53",x"27",x"03",x"BD",x"B4",x"2E",x"10",x"DE",x"75",x"7F",x"29",x"53",x"9E",x"C7",x"BF",x"2C",
    x"3E",x"8C",x"DB",x"2F",x"10",x"27",x"29",x"98",x"9E",x"38",x"BF",x"2C",x"2C",x"96",x"1A",x"B7",
    x"2C",x"2E",x"FE",x"2C",x"2A",x"30",x"41",x"27",x"1F",x"FF",x"2C",x"27",x"9E",x"38",x"9F",x"36",
    x"BE",x"2C",x"2F",x"27",x"13",x"B6",x"2C",x"29",x"26",x"0E",x"73",x"2C",x"29",x"B6",x"2C",x"31",
    x"97",x"1A",x"BD",x"DC",x"19",x"7E",x"D0",x"1A",x"BD",x"C2",x"D3",x"BD",x"D9",x"A6",x"BD",x"D9",
    x"A3",x"B6",x"2C",x"26",x"8E",x"23",x"2F",x"CE",x"D3",x"FD",x"BD",x"B0",x"02",x"BD",x"27",x"D9",
    x"BD",x"C3",x"4E",x"96",x"31",x"4C",x"27",x"03",x"BD",x"C4",x"53",x"0F",x"77",x"BD",x"C2",x"D3",
    x"BD",x"C3",x"53",x"4F",x"4B",x"0D",x"0A",x"00",x"BD",x"C6",x"63",x"BD",x"E0",x"76",x"25",x"F8",
    x"9F",x"C7",x"9D",x"C0",x"27",x"15",x"8E",x"FF",x"FF",x"9F",x"31",x"25",x"0C",x"96",x"77",x"10",
    x"26",x"FF",x"42",x"BD",x"CE",x"FB",x"7E",x"D0",x"45",x"8D",x"07",x"0D",x"78",x"27",x"D9",x"7E",
    x"D5",x"DB",x"BD",x"B7",x"8E",x"BD",x"D2",x"09",x"9E",x"33",x"BF",x"2C",x"40",x"BF",x"29",x"58",
    x"7F",x"29",x"5A",x"9E",x"C7",x"A6",x"82",x"81",x"20",x"27",x"FA",x"81",x"09",x"27",x"F6",x"A6",
    x"01",x"81",x"20",x"26",x"02",x"30",x"01",x"BD",x"CE",x"F8",x"34",x"06",x"BD",x"B3",x"E6",x"25",
    x"13",x"34",x"12",x"9F",x"6B",x"97",x"6D",x"97",x"70",x"EC",x"84",x"30",x"8B",x"9F",x"6E",x"BD",
    x"C5",x"AC",x"35",x"12",x"97",x"70",x"B6",x"29",x"5A",x"27",x"2A",x"EC",x"E4",x"31",x"8B",x"34",
    x"30",x"8D",x"24",x"35",x"50",x"11",x"83",x"9F",x"FC",x"25",x"0C",x"BD",x"D5",x"F3",x"63",x"84",
    x"8E",x"60",x"01",x"0C",x"70",x"20",x"E4",x"10",x"8E",x"29",x"56",x"35",x"06",x"ED",x"A4",x"34",
    x"20",x"31",x"AB",x"8D",x"6A",x"35",x"C0",x"10",x"AE",x"62",x"EE",x"64",x"96",x"70",x"BD",x"DC",
    x"19",x"91",x"21",x"23",x"06",x"8E",x"60",x"00",x"BD",x"D5",x"F3",x"8C",x"31",x"AB",x"EC",x"A4",
    x"27",x"31",x"33",x"CB",x"11",x"83",x"9F",x"FC",x"25",x"F2",x"34",x"20",x"31",x"AB",x"EC",x"A4",
    x"26",x"FA",x"1F",x"20",x"A3",x"E4",x"34",x"20",x"8E",x"60",x"01",x"31",x"8B",x"34",x"30",x"0C",
    x"70",x"8D",x"C4",x"35",x"70",x"96",x"70",x"97",x"6D",x"0A",x"70",x"10",x"AE",x"E4",x"BD",x"DC",
    x"32",x"35",x"20",x"EC",x"64",x"A3",x"62",x"30",x"AB",x"96",x"70",x"BD",x"DC",x"19",x"BD",x"D5",
    x"F3",x"63",x"84",x"91",x"21",x"25",x"04",x"6F",x"84",x"8D",x"0E",x"33",x"1E",x"20",x"04",x"A6",
    x"A2",x"A7",x"C2",x"10",x"AC",x"62",x"26",x"F7",x"39",x"91",x"27",x"2B",x"09",x"26",x"04",x"9C",
    x"25",x"25",x"03",x"7E",x"B1",x"FC",x"34",x"56",x"8E",x"2B",x"34",x"8D",x"07",x"35",x"56",x"97",
    x"21",x"9F",x"1F",x"39",x"CE",x"2B",x"69",x"BD",x"DC",x"09",x"73",x"2B",x"3C",x"39",x"BD",x"B6",
    x"14",x"9F",x"25",x"97",x"27",x"39",x"4F",x"8E",x"60",x"01",x"4C",x"DE",x"33",x"11",x"B3",x"2B",
    x"3C",x"26",x"06",x"BE",x"2B",x"3E",x"B6",x"2B",x"40",x"34",x"02",x"BD",x"DC",x"19",x"EC",x"84",
    x"27",x"09",x"11",x"A3",x"02",x"23",x"0D",x"30",x"8B",x"20",x"F3",x"A6",x"02",x"35",x"02",x"26",
    x"D6",x"1A",x"01",x"39",x"35",x"02",x"FF",x"2B",x"3C",x"BF",x"2B",x"3E",x"B7",x"2B",x"40",x"39",
    x"8E",x"60",x"00",x"9F",x"C7",x"86",x"01",x"97",x"1A",x"7E",x"DC",x"19",x"26",x"F1",x"8D",x"F0",
    x"4F",x"5F",x"ED",x"81",x"ED",x"81",x"4C",x"8D",x"8D",x"0F",x"72",x"0F",x"79",x"8D",x"E1",x"BD",
    x"27",x"E2",x"BD",x"D9",x"E8",x"BE",x"2C",x"4B",x"F6",x"2C",x"17",x"BD",x"B5",x"F4",x"9F",x"28",
    x"BF",x"20",x"70",x"BE",x"2D",x"17",x"B6",x"2D",x"19",x"26",x"30",x"CE",x"EF",x"81",x"BD",x"B0",
    x"02",x"BD",x"B5",x"51",x"9E",x"2E",x"96",x"30",x"10",x"BE",x"22",x"AE",x"F6",x"2C",x"4D",x"27",
    x"0C",x"BD",x"B6",x"3F",x"AF",x"A4",x"A7",x"22",x"31",x"28",x"5A",x"26",x"F4",x"BF",x"2D",x"17",
    x"B7",x"2D",x"19",x"6F",x"A4",x"CE",x"EF",x"50",x"BD",x"B0",x"02",x"DE",x"17",x"BD",x"B6",x"1F",
    x"9F",x"22",x"97",x"24",x"BF",x"2B",x"D0",x"B7",x"2B",x"D2",x"BD",x"B3",x"E1",x"C6",x"7F",x"BD",
    x"E3",x"D1",x"4F",x"5F",x"DD",x"2C",x"DD",x"2A",x"7F",x"2C",x"3E",x"DD",x"A1",x"DD",x"A3",x"F7",
    x"2C",x"29",x"FD",x"2C",x"2F",x"8D",x"4A",x"9E",x"1B",x"9F",x"1D",x"8E",x"2B",x"6A",x"33",x"88",
    x"19",x"86",x"04",x"BD",x"DC",x"0A",x"8E",x"2A",x"5E",x"BD",x"B3",x"D4",x"73",x"2B",x"15",x"8E",
    x"80",x"4F",x"BF",x"22",x"8A",x"8E",x"C7",x"52",x"BF",x"22",x"8C",x"CE",x"DF",x"7F",x"BD",x"B0",
    x"02",x"AE",x"E4",x"10",x"DE",x"28",x"6F",x"E2",x"10",x"DF",x"75",x"0F",x"36",x"0F",x"37",x"7F",
    x"29",x"53",x"6E",x"84",x"27",x"0B",x"BD",x"B7",x"8E",x"BD",x"B3",x"E6",x"24",x"08",x"7E",x"B6",
    x"D2",x"8E",x"60",x"01",x"86",x"01",x"30",x"1F",x"9F",x"3E",x"97",x"40",x"7E",x"DC",x"23",x"BD",
    x"D3",x"99",x"9D",x"C6",x"20",x"05",x"BD",x"B1",x"F2",x"1A",x"01",x"26",x"33",x"9E",x"C7",x"9F",
    x"38",x"10",x"DE",x"75",x"76",x"2B",x"D5",x"DE",x"31",x"30",x"41",x"27",x"07",x"FF",x"2C",x"27",
    x"9E",x"38",x"9F",x"36",x"8E",x"B1",x"D7",x"7D",x"2B",x"D5",x"10",x"2A",x"FD",x"5D",x"7E",x"B2",
    x"90",x"C6",x"11",x"9E",x"36",x"26",x"02",x"0E",x"B7",x"9F",x"C7",x"BE",x"2C",x"27",x"9F",x"31",
    x"39",x"CE",x"EF",x"A2",x"7E",x"B0",x"02",x"F6",x"2C",x"4D",x"34",x"04",x"B6",x"2C",x"17",x"D6",
    x"30",x"9E",x"2E",x"10",x"9E",x"17",x"FE",x"2C",x"4B",x"34",x"76",x"9D",x"C6",x"27",x"43",x"81",
    x"2C",x"27",x"05",x"BD",x"C1",x"66",x"AF",x"64",x"BD",x"B8",x"E7",x"27",x"1A",x"96",x"4D",x"A7",
    x"61",x"BD",x"C1",x"66",x"8C",x"9F",x"FF",x"22",x"6E",x"8C",x"60",x"00",x"24",x"07",x"AF",x"66",
    x"8D",x"60",x"8E",x"60",x"00",x"AF",x"62",x"BD",x"B8",x"E7",x"27",x"0B",x"C6",x"80",x"BD",x"C1",
    x"E9",x"E7",x"E4",x"AE",x"66",x"8D",x"4D",x"9D",x"C6",x"27",x"07",x"BD",x"C1",x"64",x"AF",x"66",
    x"8D",x"40",x"A6",x"61",x"AE",x"62",x"8D",x"5C",x"8D",x"97",x"E6",x"68",x"27",x"05",x"8D",x"7F",
    x"5A",x"26",x"FB",x"8D",x"4F",x"EE",x"64",x"8D",x"56",x"8D",x"49",x"35",x"36",x"B7",x"2C",x"17",
    x"D7",x"30",x"9F",x"2E",x"10",x"9F",x"17",x"35",x"10",x"BF",x"2C",x"4B",x"35",x"44",x"F7",x"2C",
    x"4D",x"F6",x"2C",x"17",x"8D",x"0E",x"9F",x"28",x"1F",x"14",x"34",x"40",x"7F",x"2D",x"19",x"7E",
    x"B4",x"3F",x"E6",x"62",x"8C",x"5F",x"FF",x"22",x"18",x"86",x"08",x"3D",x"40",x"50",x"82",x"00",
    x"30",x"8B",x"34",x"10",x"1F",x"10",x"83",x"00",x"5A",x"23",x"06",x"93",x"1B",x"23",x"02",x"35",
    x"90",x"7E",x"B1",x"FC",x"91",x"21",x"2B",x"F9",x"26",x"04",x"9C",x"1F",x"23",x"F3",x"39",x"34",
    x"12",x"1F",x"30",x"20",x"04",x"6A",x"E4",x"80",x"40",x"81",x"40",x"24",x"F8",x"34",x"06",x"EC",
    x"63",x"A3",x"E1",x"81",x"60",x"24",x"04",x"6A",x"E4",x"8B",x"40",x"ED",x"61",x"35",x"92",x"34",
    x"46",x"1F",x"10",x"A3",x"62",x"81",x"60",x"24",x"07",x"6A",x"E4",x"CC",x"9F",x"FF",x"A3",x"62",
    x"1F",x"01",x"35",x"C6",x"81",x"22",x"10",x"27",x"1E",x"37",x"BD",x"D3",x"99",x"9D",x"C6",x"10",
    x"27",x"FD",x"DA",x"BD",x"B4",x"3F",x"20",x"1B",x"1F",x"89",x"9D",x"C0",x"C1",x"BB",x"27",x"18",
    x"C1",x"BC",x"26",x"62",x"C6",x"03",x"BD",x"B1",x"E1",x"DE",x"C7",x"9E",x"31",x"86",x"BC",x"D6",
    x"1A",x"34",x"56",x"8D",x"03",x"7E",x"D0",x"05",x"9D",x"C6",x"BD",x"B7",x"8E",x"8D",x"60",x"30",
    x"01",x"DC",x"33",x"10",x"93",x"31",x"22",x"05",x"BD",x"B3",x"E6",x"20",x"05",x"96",x"1A",x"BD",
    x"B3",x"EB",x"25",x"2E",x"97",x"1A",x"30",x"1F",x"9F",x"C7",x"39",x"BE",x"2C",x"3C",x"9F",x"33",
    x"30",x"01",x"26",x"E4",x"32",x"62",x"7E",x"B2",x"9B",x"26",x"EF",x"86",x"FF",x"97",x"48",x"86",
    x"81",x"BD",x"E4",x"A2",x"32",x"84",x"9F",x"75",x"81",x"BC",x"27",x"0D",x"BD",x"28",x"09",x"C6",
    x"03",x"8C",x"C6",x"08",x"0E",x"B7",x"7E",x"B8",x"F4",x"35",x"56",x"9F",x"31",x"DF",x"C7",x"D7",
    x"1A",x"BD",x"DC",x"23",x"8D",x"06",x"8C",x"8D",x"06",x"9F",x"C7",x"39",x"C6",x"3A",x"86",x"5F",
    x"9E",x"C7",x"D7",x"00",x"5F",x"1F",x"98",x"D6",x"00",x"97",x"00",x"A6",x"84",x"27",x"EC",x"34",
    x"04",x"A1",x"E0",x"27",x"E6",x"30",x"01",x"81",x"22",x"27",x"EA",x"4C",x"26",x"02",x"30",x"01",
    x"81",x"8A",x"26",x"E7",x"0C",x"66",x"20",x"E3",x"BD",x"B9",x"06",x"9D",x"C6",x"81",x"87",x"26",
    x"0C",x"9E",x"C7",x"9D",x"C0",x"9F",x"C7",x"81",x"BB",x"27",x"06",x"20",x"A9",x"C6",x"C4",x"9D",
    x"BD",x"CE",x"C2",x"56",x"BD",x"B0",x"02",x"5D",x"26",x"13",x"0F",x"66",x"8D",x"A6",x"4D",x"27",
    x"AA",x"9D",x"C0",x"81",x"8F",x"26",x"F5",x"0A",x"66",x"2A",x"F1",x"9D",x"C0",x"9D",x"C6",x"10",
    x"25",x"FF",x"35",x"7E",x"D0",x"4B",x"81",x"98",x"10",x"27",x"11",x"34",x"81",x"B0",x"10",x"27",
    x"12",x"6B",x"81",x"AF",x"10",x"27",x"12",x"4E",x"BD",x"C1",x"4E",x"C6",x"87",x"9D",x"BD",x"34",
    x"02",x"81",x"BC",x"27",x"04",x"81",x"BB",x"26",x"B2",x"0A",x"51",x"26",x"05",x"35",x"04",x"7E",
    x"B6",x"6A",x"9D",x"C0",x"8D",x"08",x"81",x"2C",x"27",x"EF",x"9D",x"C6",x"35",x"84",x"8E",x"00",
    x"00",x"9F",x"33",x"25",x"02",x"0E",x"C6",x"80",x"30",x"97",x"00",x"DC",x"33",x"81",x"18",x"22",
    x"8A",x"58",x"49",x"58",x"49",x"D3",x"33",x"58",x"49",x"DB",x"00",x"89",x"00",x"DD",x"33",x"9D",
    x"C0",x"20",x"E0",x"BD",x"BB",x"96",x"9F",x"48",x"97",x"4A",x"8D",x"45",x"C6",x"D4",x"9D",x"BD",
    x"96",x"05",x"34",x"02",x"BD",x"B9",x"06",x"35",x"02",x"BD",x"B0",x"27",x"7E",x"B9",x"45",x"8D",
    x"E2",x"27",x"05",x"BD",x"B0",x"2C",x"20",x"29",x"DE",x"48",x"96",x"4A",x"BD",x"DC",x"27",x"AE",
    x"41",x"9C",x"17",x"25",x"06",x"C6",x"44",x"6D",x"C4",x"26",x"1B",x"D6",x"51",x"E1",x"C4",x"23",
    x"0B",x"34",x"40",x"6F",x"C4",x"BD",x"BF",x"C0",x"35",x"40",x"AF",x"41",x"E7",x"C4",x"BD",x"BE",
    x"37",x"7E",x"DC",x"23",x"C6",x"16",x"0E",x"B7",x"BD",x"27",x"D3",x"9D",x"C0",x"27",x"F5",x"24",
    x"0C",x"10",x"9E",x"C7",x"CE",x"C4",x"0A",x"8D",x"37",x"10",x"9F",x"C7",x"39",x"81",x"41",x"2D",
    x"1B",x"BD",x"BB",x"7C",x"BD",x"B9",x"45",x"26",x"0B",x"E6",x"84",x"D7",x"51",x"AE",x"01",x"BD",
    x"BE",x"1E",x"20",x"05",x"CE",x"C1",x"84",x"8D",x"17",x"7E",x"DC",x"23",x"81",x"2E",x"27",x"D1",
    x"81",x"26",x"27",x"CD",x"81",x"C8",x"26",x"0B",x"86",x"7D",x"BD",x"B9",x"0C",x"CE",x"CC",x"44",
    x"7E",x"B0",x"02",x"81",x"C7",x"27",x"B1",x"81",x"22",x"26",x"08",x"9E",x"C7",x"BD",x"BF",x"90",
    x"9F",x"C7",x"39",x"81",x"C5",x"26",x"0D",x"86",x"5A",x"BD",x"B9",x"0C",x"BD",x"B0",x"22",x"03",
    x"50",x"03",x"51",x"39",x"81",x"C2",x"26",x"08",x"F6",x"2C",x"26",x"9D",x"C0",x"7E",x"BD",x"D6",
    x"81",x"C1",x"26",x"0D",x"9D",x"C0",x"BE",x"2C",x"2A",x"9F",x"50",x"CE",x"CB",x"A9",x"7E",x"B0",
    x"02",x"81",x"C0",x"10",x"27",x"10",x"C3",x"81",x"BD",x"10",x"27",x"34",x"99",x"4C",x"26",x"33",
    x"9D",x"C0",x"1F",x"89",x"58",x"9D",x"C0",x"C1",x"80",x"23",x"04",x"6E",x"9F",x"27",x"82",x"BE",
    x"27",x"78",x"3A",x"AE",x"84",x"2A",x"0D",x"30",x"89",x"30",x"00",x"34",x"10",x"8D",x"14",x"35",
    x"40",x"7E",x"B0",x"02",x"8C",x"40",x"00",x"25",x"04",x"6E",x"89",x"70",x"00",x"30",x"89",x"B0",
    x"00",x"34",x"10",x"8D",x"05",x"8D",x"2F",x"C6",x"29",x"8C",x"C6",x"28",x"8C",x"C6",x"2C",x"E1",
    x"9F",x"21",x"C7",x"26",x"0F",x"0E",x"C0",x"9D",x"C6",x"27",x"08",x"81",x"2C",x"26",x"05",x"9D",
    x"C0",x"81",x"2C",x"39",x"C6",x"02",x"0E",x"B7",x"8D",x"0C",x"8D",x"49",x"26",x"4B",x"7E",x"BF",
    x"3D",x"9E",x"C7",x"7E",x"B6",x"A6",x"8D",x"F9",x"4F",x"8C",x"96",x"4B",x"34",x"02",x"C6",x"01",
    x"BD",x"B1",x"E1",x"BD",x"B8",x"08",x"0F",x"03",x"6F",x"E2",x"9E",x"C7",x"BF",x"2C",x"32",x"9D",
    x"C6",x"80",x"D3",x"25",x"13",x"81",x"03",x"24",x"0F",x"81",x"01",x"49",x"A8",x"E4",x"A1",x"E4",
    x"25",x"C2",x"A7",x"E4",x"9D",x"C0",x"20",x"E9",x"E6",x"E0",x"10",x"26",x"00",x"F8",x"25",x"0A",
    x"35",x"82",x"86",x"04",x"8C",x"86",x"03",x"90",x"05",x"39",x"8B",x"0C",x"24",x"F2",x"1F",x"89",
    x"26",x"06",x"8D",x"F1",x"10",x"27",x"05",x"AC",x"34",x"04",x"58",x"EB",x"E0",x"8E",x"B0",x"BF",
    x"3A",x"A6",x"E4",x"E6",x"84",x"A1",x"84",x"24",x"D7",x"8D",x"8F",x"8D",x"02",x"20",x"A7",x"D7",
    x"4B",x"10",x"8E",x"B8",x"BF",x"EE",x"01",x"34",x"60",x"C1",x"51",x"25",x"6A",x"C4",x"FE",x"C1",
    x"7A",x"27",x"64",x"8D",x"70",x"8D",x"83",x"BD",x"B8",x"FA",x"BD",x"BA",x"16",x"D6",x"4C",x"D1",
    x"05",x"27",x"0C",x"C1",x"08",x"26",x"0D",x"CE",x"CB",x"5A",x"8D",x"48",x"0C",x"03",x"39",x"C1",
    x"08",x"27",x"F9",x"39",x"8D",x"9C",x"24",x"2F",x"D7",x"05",x"8D",x"02",x"8D",x"E9",x"DC",x"5F",
    x"9E",x"54",x"9F",x"5F",x"DD",x"54",x"DC",x"5D",x"9E",x"52",x"9F",x"5D",x"DD",x"52",x"DC",x"59",
    x"9E",x"4E",x"9F",x"59",x"DD",x"4E",x"96",x"61",x"D6",x"56",x"D7",x"61",x"97",x"56",x"DC",x"5B",
    x"9E",x"50",x"9F",x"5B",x"DD",x"50",x"39",x"26",x"08",x"D7",x"05",x"8D",x"E1",x"8D",x"02",x"20",
    x"DD",x"CE",x"CB",x"6D",x"7E",x"B0",x"02",x"BD",x"B0",x"22",x"8D",x"09",x"BD",x"B9",x"0A",x"BD",
    x"B0",x"22",x"8D",x"22",x"39",x"35",x"20",x"CE",x"21",x"52",x"D6",x"05",x"C1",x"04",x"23",x"02",
    x"33",x"44",x"25",x"04",x"96",x"56",x"34",x"02",x"54",x"AE",x"C3",x"34",x"10",x"5A",x"26",x"F9",
    x"D6",x"05",x"34",x"04",x"6E",x"A4",x"35",x"20",x"35",x"14",x"D7",x"4C",x"C1",x"02",x"27",x"12",
    x"CE",x"21",x"59",x"8C",x"35",x"10",x"AF",x"C1",x"C0",x"02",x"26",x"F8",x"35",x"04",x"D7",x"61",
    x"6E",x"A4",x"9F",x"5B",x"6E",x"A4",x"A6",x"E4",x"81",x"64",x"25",x"07",x"BE",x"2C",x"32",x"9F",
    x"C7",x"35",x"82",x"BD",x"B9",x"01",x"34",x"04",x"8D",x"0F",x"CB",x"01",x"59",x"E4",x"E0",x"27",
    x"02",x"C6",x"FF",x"BD",x"BD",x"D4",x"7E",x"B9",x"16",x"C6",x"64",x"BD",x"B9",x"45",x"27",x"06",
    x"8E",x"B0",x"E2",x"7E",x"B9",x"6F",x"BD",x"BF",x"4A",x"86",x"64",x"BD",x"B9",x"0C",x"BD",x"BF",
    x"38",x"BD",x"BE",x"75",x"A6",x"E4",x"90",x"51",x"27",x"07",x"86",x"FF",x"24",x"03",x"E6",x"E4",
    x"40",x"97",x"56",x"30",x"61",x"5C",x"5A",x"26",x"04",x"D6",x"56",x"20",x"0D",x"A6",x"80",x"A1",
    x"C0",x"27",x"F3",x"C6",x"FF",x"24",x"01",x"50",x"D7",x"56",x"BD",x"BE",x"CB",x"D6",x"56",x"39",
    x"9D",x"BA",x"BD",x"B9",x"06",x"BD",x"B0",x"22",x"9E",x"50",x"39",x"9D",x"BA",x"BD",x"B9",x"06",
    x"CE",x"CB",x"6D",x"BD",x"B0",x"02",x"8E",x"21",x"4E",x"39",x"04",x"00",x"08",x"03",x"02",x"CE",
    x"2B",x"84",x"9E",x"C7",x"A6",x"84",x"5F",x"20",x"08",x"30",x"01",x"A6",x"84",x"9D",x"CD",x"25",
    x"08",x"81",x"41",x"25",x"0D",x"81",x"5A",x"22",x"09",x"C1",x"10",x"27",x"EC",x"A7",x"C0",x"5C",
    x"20",x"E7",x"D7",x"44",x"10",x"27",x"FE",x"0C",x"CE",x"BA",x"BA",x"80",x"21",x"81",x"04",x"23",
    x"08",x"CE",x"2B",x"29",x"B6",x"2B",x"84",x"30",x"1F",x"E6",x"C6",x"27",x"F4",x"DA",x"04",x"9F",
    x"C7",x"9D",x"C0",x"0D",x"04",x"26",x"06",x"81",x"28",x"26",x"02",x"CA",x"80",x"D7",x"05",x"39",
    x"0F",x"04",x"BD",x"28",x"00",x"8D",x"A8",x"D6",x"44",x"5A",x"26",x"1B",x"96",x"05",x"81",x"03",
    x"27",x"15",x"81",x"04",x"22",x"11",x"8E",x"2A",x"5D",x"B6",x"2B",x"84",x"80",x"41",x"C6",x"07",
    x"3D",x"DB",x"05",x"3A",x"1A",x"01",x"39",x"DC",x"1B",x"83",x"00",x"04",x"DD",x"D6",x"DE",x"1D",
    x"DF",x"D8",x"DC",x"D6",x"D3",x"D8",x"46",x"56",x"C4",x"FC",x"1F",x"03",x"A6",x"43",x"91",x"05",
    x"26",x"1F",x"A6",x"42",x"BD",x"DC",x"27",x"AE",x"C4",x"E6",x"80",x"D1",x"44",x"26",x"12",x"10",
    x"8E",x"2B",x"84",x"A6",x"80",x"A1",x"A0",x"26",x"08",x"5A",x"26",x"F7",x"96",x"8B",x"1C",x"FE",
    x"39",x"24",x"CD",x"11",x"93",x"D6",x"27",x"F6",x"DF",x"D6",x"20",x"C6",x"8D",x"92",x"26",x"1F",
    x"0D",x"05",x"2A",x"0D",x"BD",x"BD",x"5A",x"8E",x"00",x"0A",x"AC",x"E1",x"25",x"26",x"5A",x"26",
    x"F9",x"8E",x"2D",x"1B",x"20",x"33",x"9E",x"C7",x"9F",x"3A",x"BD",x"BB",x"10",x"27",x"19",x"25",
    x"30",x"0D",x"05",x"2A",x"24",x"BD",x"BD",x"5A",x"E1",x"80",x"26",x"08",x"BD",x"BC",x"C1",x"BD",
    x"DC",x"19",x"20",x"15",x"C6",x"09",x"0E",x"B7",x"D6",x"05",x"2B",x"1A",x"5C",x"DB",x"44",x"8D",
    x"2E",x"8D",x"3D",x"8D",x"1B",x"6F",x"84",x"6F",x"01",x"96",x"05",x"84",x"0F",x"97",x"05",x"96",
    x"8B",x"9F",x"45",x"97",x"47",x"39",x"0F",x"06",x"8D",x"5A",x"9E",x"3A",x"9F",x"C7",x"20",x"B6",
    x"CE",x"2B",x"84",x"D6",x"44",x"E7",x"80",x"A6",x"C0",x"A7",x"80",x"5A",x"26",x"F9",x"39",x"4F",
    x"34",x"46",x"1F",x"03",x"9E",x"25",x"96",x"27",x"BD",x"B6",x"3F",x"BD",x"B3",x"DE",x"35",x"C6",
    x"C6",x"02",x"BD",x"B1",x"E1",x"33",x"44",x"34",x"40",x"10",x"9E",x"1D",x"33",x"24",x"DF",x"1D",
    x"BD",x"B3",x"B3",x"35",x"40",x"96",x"27",x"BD",x"DC",x"19",x"9E",x"25",x"AF",x"C4",x"96",x"8B",
    x"D6",x"05",x"ED",x"42",x"39",x"C6",x"80",x"D7",x"04",x"D7",x"06",x"BD",x"BB",x"12",x"27",x"04",
    x"C6",x"0A",x"0E",x"B7",x"FF",x"2B",x"A5",x"8E",x"2B",x"94",x"8D",x"A4",x"BD",x"BD",x"5A",x"58",
    x"CB",x"07",x"FB",x"2B",x"94",x"8D",x"A8",x"96",x"26",x"84",x"FE",x"97",x"26",x"FE",x"2B",x"A5",
    x"8D",x"AE",x"9F",x"45",x"96",x"27",x"97",x"47",x"CE",x"2B",x"94",x"E6",x"C0",x"6F",x"80",x"8D",
    x"86",x"D6",x"DA",x"E7",x"80",x"1F",x"42",x"34",x"10",x"EE",x"A4",x"0D",x"06",x"26",x"03",x"CE",
    x"00",x"0A",x"EF",x"A1",x"33",x"41",x"EF",x"81",x"5A",x"26",x"EE",x"DE",x"45",x"EF",x"81",x"96",
    x"47",x"A7",x"80",x"9F",x"0A",x"35",x"10",x"8D",x"37",x"DE",x"DD",x"EF",x"9F",x"21",x"0A",x"BD",
    x"B3",x"DE",x"20",x"0B",x"6F",x"80",x"8C",x"A0",x"00",x"26",x"F9",x"4C",x"8E",x"60",x"00",x"BD",
    x"DC",x"19",x"91",x"47",x"26",x"EE",x"6F",x"80",x"9C",x"45",x"26",x"FA",x"F6",x"2B",x"94",x"E7",
    x"84",x"7E",x"DC",x"23",x"9D",x"C0",x"BD",x"BC",x"25",x"9D",x"C6",x"81",x"2C",x"27",x"F5",x"39",
    x"86",x"4F",x"97",x"04",x"96",x"05",x"84",x"0F",x"97",x"05",x"4F",x"5F",x"DD",x"DB",x"5C",x"DD",
    x"DD",x"35",x"20",x"EC",x"E1",x"34",x"20",x"8D",x"3A",x"0A",x"DA",x"26",x"F4",x"DC",x"DB",x"C3",
    x"00",x"01",x"DD",x"DD",x"4F",x"D6",x"05",x"8D",x"3E",x"6F",x"E2",x"20",x"05",x"83",x"3F",x"F8",
    x"6C",x"E4",x"10",x"83",x"3F",x"F8",x"24",x"F5",x"34",x"06",x"EC",x"81",x"A3",x"E1",x"81",x"60",
    x"24",x"05",x"C3",x"3F",x"F8",x"6C",x"E4",x"DD",x"DB",x"A6",x"84",x"A0",x"E0",x"9E",x"DB",x"39",
    x"7E",x"BB",x"B4",x"10",x"A3",x"84",x"24",x"F8",x"8D",x"0D",x"D3",x"DB",x"2B",x"F2",x"DD",x"DB",
    x"EC",x"81",x"8D",x"03",x"DD",x"DD",x"39",x"DE",x"DD",x"91",x"DD",x"23",x"02",x"1E",x"03",x"4D",
    x"26",x"DE",x"D7",x"4F",x"DF",x"50",x"96",x"51",x"3D",x"34",x"06",x"DC",x"4F",x"3D",x"4D",x"26",
    x"CF",x"EB",x"E4",x"E7",x"E4",x"25",x"C9",x"35",x"86",x"9D",x"C0",x"BD",x"B8",x"F8",x"BD",x"B0",
    x"22",x"9E",x"50",x"DC",x"50",x"2A",x"CF",x"7E",x"BF",x"43",x"35",x"20",x"96",x"8B",x"D6",x"05",
    x"1F",x"03",x"BD",x"DC",x"23",x"0F",x"DA",x"96",x"DA",x"34",x"72",x"8D",x"DC",x"35",x"72",x"4C",
    x"97",x"DA",x"2B",x"E3",x"DC",x"50",x"34",x"06",x"9D",x"C6",x"81",x"2C",x"27",x"E9",x"BD",x"B8",
    x"D7",x"1F",x"30",x"BD",x"DC",x"27",x"D7",x"05",x"D6",x"DA",x"6E",x"A4",x"BD",x"BB",x"96",x"D6",
    x"05",x"34",x"16",x"8D",x"27",x"9D",x"BA",x"BD",x"BB",x"96",x"D6",x"05",x"E1",x"61",x"10",x"26",
    x"01",x"9B",x"9F",x"45",x"97",x"47",x"CE",x"21",x"4E",x"BD",x"DC",x"01",x"35",x"16",x"BD",x"DC",
    x"27",x"8D",x"0C",x"9E",x"45",x"96",x"47",x"BD",x"DC",x"27",x"8D",x"03",x"7E",x"DC",x"23",x"CE",
    x"21",x"4E",x"D6",x"05",x"34",x"04",x"A6",x"84",x"E6",x"C4",x"A7",x"C0",x"E7",x"80",x"6A",x"E4",
    x"26",x"F4",x"35",x"84",x"1D",x"21",x"4F",x"DD",x"50",x"86",x"02",x"97",x"05",x"39",x"C6",x"01",
    x"9D",x"C6",x"81",x"28",x"26",x"04",x"BD",x"B8",x"D3",x"8C",x"8D",x"EA",x"CE",x"CA",x"B8",x"7E",
    x"B0",x"02",x"CE",x"CF",x"6D",x"20",x"03",x"CE",x"CF",x"5D",x"34",x"40",x"BD",x"B8",x"F8",x"9D",
    x"C6",x"81",x"2C",x"27",x"05",x"35",x"40",x"7E",x"B8",x"D7",x"BD",x"B9",x"F5",x"9D",x"C0",x"BD",
    x"B8",x"F8",x"BD",x"BA",x"16",x"BD",x"B9",x"8D",x"EE",x"E4",x"8D",x"D3",x"20",x"E1",x"8D",x"0B",
    x"23",x"1B",x"A6",x"80",x"A7",x"C0",x"8D",x"53",x"26",x"F8",x"39",x"8D",x"1C",x"27",x"06",x"34",
    x"10",x"3A",x"8C",x"9F",x"FF",x"35",x"90",x"8D",x"F2",x"22",x"05",x"1E",x"13",x"7E",x"DC",x"01",
    x"A6",x"C0",x"A7",x"80",x"8D",x"35",x"26",x"F8",x"39",x"9C",x"17",x"25",x"0A",x"1F",x"10",x"93",
    x"17",x"9E",x"87",x"30",x"8B",x"20",x"1E",x"96",x"24",x"97",x"50",x"1F",x"10",x"20",x"04",x"80",
    x"40",x"0C",x"50",x"81",x"40",x"24",x"F8",x"D3",x"22",x"81",x"A0",x"25",x"04",x"80",x"40",x"0C",
    x"50",x"1F",x"01",x"8D",x"13",x"CE",x"23",x"2F",x"D6",x"51",x"39",x"5A",x"27",x"CA",x"8C",x"A0",
    x"00",x"26",x"C5",x"0C",x"50",x"8E",x"60",x"00",x"96",x"50",x"7E",x"DC",x"19",x"BD",x"B8",x"DA",
    x"BD",x"BF",x"30",x"35",x"10",x"BD",x"BF",x"4A",x"34",x"10",x"7E",x"C1",x"60",x"8D",x"EE",x"4F",
    x"20",x"20",x"8D",x"E9",x"5D",x"27",x"53",x"5A",x"34",x"04",x"C6",x"FF",x"9D",x"C6",x"81",x"29",
    x"27",x"03",x"BD",x"C1",x"60",x"35",x"02",x"20",x"09",x"8D",x"D2",x"1F",x"98",x"A0",x"E4",x"24",
    x"DE",x"40",x"8D",x"08",x"7E",x"B8",x"D7",x"4F",x"E6",x"62",x"21",x"5F",x"35",x"20",x"DD",x"50",
    x"35",x"04",x"30",x"E4",x"3A",x"34",x"10",x"D6",x"50",x"30",x"62",x"3A",x"8D",x"97",x"27",x"0E",
    x"AC",x"E4",x"24",x"07",x"A6",x"80",x"A7",x"C0",x"5A",x"26",x"F5",x"D0",x"51",x"50",x"10",x"EE",
    x"E4",x"34",x"20",x"20",x"73",x"8D",x"41",x"17",x"FF",x"7B",x"27",x"47",x"E6",x"C4",x"39",x"8D",
    x"F4",x"7E",x"BD",x"D6",x"8D",x"44",x"BD",x"B8",x"08",x"8D",x"2D",x"BD",x"BE",x"75",x"EB",x"E4",
    x"25",x"2E",x"D7",x"4F",x"1F",x"31",x"4F",x"33",x"CB",x"D6",x"51",x"27",x"08",x"3A",x"A6",x"82",
    x"A7",x"C2",x"5A",x"26",x"F9",x"8D",x"A0",x"D6",x"4F",x"8D",x"3D",x"7E",x"B9",x"16",x"9D",x"BA",
    x"BD",x"B9",x"06",x"8E",x"23",x"2F",x"D6",x"51",x"BD",x"B9",x"45",x"27",x"31",x"C6",x"0D",x"8C",
    x"C6",x"0F",x"8C",x"C6",x"05",x"8C",x"C6",x"0E",x"0E",x"B7",x"35",x"20",x"BD",x"BE",x"75",x"4F",
    x"34",x"06",x"BD",x"B1",x"E3",x"EC",x"E1",x"27",x"0B",x"33",x"CB",x"A6",x"C2",x"34",x"02",x"5A",
    x"26",x"F9",x"D6",x"51",x"34",x"04",x"6E",x"A4",x"D7",x"51",x"86",x"03",x"97",x"05",x"39",x"86",
    x"4F",x"34",x"02",x"BD",x"C1",x"69",x"35",x"02",x"CE",x"C4",x"D4",x"8D",x"05",x"20",x"0F",x"CE",
    x"C5",x"16",x"10",x"8E",x"2B",x"A7",x"7E",x"B0",x"02",x"BD",x"B8",x"FA",x"8D",x"F1",x"30",x"1F",
    x"86",x"22",x"1F",x"89",x"30",x"01",x"DD",x"00",x"5F",x"CE",x"23",x"2F",x"A6",x"80",x"27",x"0D",
    x"91",x"00",x"27",x"09",x"91",x"01",x"27",x"05",x"A7",x"C0",x"5C",x"20",x"EF",x"81",x"22",x"27",
    x"B7",x"30",x"1F",x"20",x"B3",x"32",x"62",x"8D",x"91",x"8D",x"14",x"27",x"89",x"BD",x"BE",x"C7",
    x"D6",x"51",x"9E",x"2C",x"34",x"10",x"3A",x"9C",x"17",x"22",x"EA",x"9F",x"2C",x"35",x"90",x"BD",
    x"28",x"03",x"0F",x"EE",x"0F",x"EF",x"DC",x"2C",x"DD",x"F0",x"DE",x"1B",x"20",x"39",x"E6",x"43",
    x"C5",x"41",x"27",x"31",x"A6",x"42",x"BD",x"DC",x"27",x"AE",x"C4",x"E6",x"80",x"3A",x"6D",x"43",
    x"2A",x"21",x"E6",x"80",x"58",x"3A",x"10",x"AE",x"03",x"A6",x"02",x"AE",x"84",x"30",x"1D",x"8C",
    x"60",x"00",x"24",x"08",x"30",x"89",x"3F",x"F8",x"4A",x"BD",x"DC",x"19",x"8D",x"59",x"31",x"3F",
    x"26",x"EB",x"8C",x"8D",x"52",x"33",x"44",x"11",x"93",x"1D",x"26",x"C2",x"CE",x"21",x"2A",x"20",
    x"04",x"30",x"42",x"8D",x"42",x"EE",x"C4",x"26",x"F8",x"86",x"0A",x"8E",x"2B",x"16",x"8D",x"37",
    x"30",x"03",x"4A",x"26",x"F9",x"BD",x"28",x"06",x"DC",x"2C",x"10",x"93",x"F0",x"27",x"21",x"DE",
    x"EB",x"96",x"ED",x"BD",x"DC",x"27",x"E6",x"C4",x"D7",x"51",x"9E",x"EE",x"AF",x"41",x"34",x"10",
    x"3A",x"9F",x"EE",x"9E",x"F0",x"BD",x"BE",x"1E",x"35",x"10",x"BD",x"BE",x"37",x"16",x"FF",x"76",
    x"9E",x"EE",x"9F",x"2C",x"93",x"EE",x"39",x"34",x"02",x"A6",x"84",x"27",x"16",x"EC",x"01",x"10",
    x"93",x"F0",x"22",x"0F",x"10",x"93",x"EE",x"25",x"0A",x"27",x"0A",x"DD",x"F0",x"96",x"8B",x"9F",
    x"EB",x"97",x"ED",x"35",x"82",x"EB",x"84",x"89",x"00",x"DD",x"EE",x"35",x"82",x"BD",x"B8",x"DA",
    x"BD",x"C1",x"4E",x"34",x"04",x"9D",x"BA",x"BD",x"E3",x"EB",x"34",x"04",x"BD",x"B8",x"D7",x"35",
    x"06",x"20",x"05",x"BD",x"C1",x"55",x"86",x"20",x"D7",x"51",x"27",x"08",x"8E",x"23",x"2F",x"A7",
    x"80",x"5A",x"26",x"FB",x"7E",x"BF",x"6A",x"86",x"4F",x"34",x"02",x"BD",x"B7",x"B3",x"10",x"26",
    x"FE",x"7B",x"9E",x"48",x"96",x"4A",x"BD",x"DC",x"27",x"BD",x"BE",x"75",x"E0",x"84",x"25",x"0E",
    x"E6",x"84",x"D7",x"51",x"AE",x"01",x"BD",x"BE",x"37",x"BD",x"DC",x"23",x"35",x"82",x"50",x"34",
    x"04",x"D6",x"51",x"4F",x"31",x"CB",x"6D",x"61",x"27",x"0F",x"E6",x"E4",x"33",x"AB",x"D6",x"51",
    x"27",x"07",x"A6",x"A2",x"A7",x"C2",x"5A",x"26",x"F9",x"35",x"04",x"86",x"20",x"A7",x"A0",x"5A",
    x"26",x"FB",x"20",x"CC",x"8D",x"1C",x"BD",x"BF",x"33",x"4F",x"A7",x"8B",x"BD",x"CF",x"05",x"83",
    x"00",x"05",x"4D",x"10",x"26",x"FE",x"29",x"D7",x"51",x"CE",x"23",x"2F",x"8E",x"29",x"5A",x"7E",
    x"DC",x"01",x"9E",x"31",x"30",x"01",x"26",x"23",x"C6",x"0C",x"0E",x"B7",x"BD",x"BF",x"33",x"9E",
    x"C7",x"34",x"10",x"6F",x"E2",x"BD",x"BF",x"4A",x"30",x"61",x"9F",x"C7",x"BD",x"B9",x"06",x"BD",
    x"C5",x"2B",x"35",x"04",x"4F",x"32",x"EB",x"35",x"12",x"9F",x"C7",x"39",x"9D",x"C0",x"BD",x"B8",
    x"F8",x"8D",x"02",x"0E",x"C6",x"BD",x"B0",x"22",x"DC",x"50",x"4D",x"10",x"26",x"FD",x"E4",x"39",
    x"9D",x"BA",x"20",x"EA",x"9D",x"BA",x"BD",x"B9",x"06",x"CE",x"CD",x"CA",x"7E",x"B0",x"02",x"81",
    x"24",x"34",x"01",x"26",x"02",x"9D",x"C0",x"BD",x"B8",x"DA",x"8D",x"EA",x"35",x"01",x"34",x"10",
    x"27",x"09",x"8D",x"5D",x"E6",x"F1",x"BD",x"BD",x"D6",x"20",x"0F",x"8D",x"D3",x"8D",x"52",x"CE",
    x"23",x"2F",x"35",x"10",x"BD",x"BF",x"68",x"BD",x"DC",x"01",x"8D",x"42",x"7E",x"B8",x"D7",x"8D",
    x"C5",x"34",x"10",x"BD",x"B9",x"08",x"8D",x"39",x"BD",x"B9",x"45",x"27",x"06",x"8D",x"A6",x"E7",
    x"F1",x"20",x"2B",x"8E",x"23",x"2F",x"35",x"40",x"D6",x"51",x"27",x"22",x"BD",x"DC",x"01",x"20",
    x"1D",x"8D",x"A3",x"34",x"10",x"8D",x"99",x"D7",x"48",x"5F",x"9D",x"C6",x"27",x"02",x"8D",x"90",
    x"D7",x"49",x"8D",x"0D",x"35",x"10",x"A6",x"84",x"98",x"49",x"94",x"48",x"27",x"F8",x"7E",x"DC",
    x"23",x"96",x"4D",x"BD",x"DC",x"19",x"7E",x"D2",x"03",x"34",x"04",x"BD",x"C1",x"4E",x"E1",x"E0",
    x"23",x"0E",x"7E",x"BF",x"43",x"D6",x"8C",x"8D",x"F0",x"5D",x"26",x"02",x"D6",x"8C",x"D7",x"4D",
    x"39",x"D6",x"4D",x"7E",x"BD",x"D6",x"27",x"06",x"BD",x"C1",x"66",x"BF",x"27",x"A8",x"8D",x"D1",
    x"FE",x"27",x"A8",x"BD",x"B0",x"0E",x"20",x"C6",x"BD",x"B9",x"45",x"27",x"09",x"BD",x"C1",x"55",
    x"CE",x"D3",x"BB",x"7E",x"B0",x"02",x"BD",x"BF",x"CF",x"BD",x"DC",x"23",x"DC",x"17",x"93",x"2C",
    x"DD",x"50",x"7E",x"B8",x"8B",x"BD",x"B9",x"08",x"BD",x"B0",x"22",x"9D",x"C6",x"81",x"29",x"10",
    x"26",x"F6",x"B1",x"DC",x"50",x"2A",x"02",x"4F",x"5F",x"DD",x"5B",x"4F",x"BD",x"D6",x"C4",x"F6",
    x"2C",x"37",x"26",x"01",x"4C",x"DD",x"50",x"CE",x"CC",x"98",x"BD",x"B0",x"02",x"D6",x"51",x"F0",
    x"2C",x"36",x"24",x"04",x"8D",x"77",x"D6",x"51",x"7E",x"C3",x"0E",x"27",x"70",x"8D",x"0B",x"0F",
    x"77",x"39",x"BD",x"D3",x"A7",x"BD",x"D6",x"F9",x"0E",x"C6",x"81",x"23",x"26",x"06",x"8D",x"F2",
    x"27",x"5B",x"9D",x"BA",x"81",x"BF",x"10",x"27",x"04",x"A0",x"26",x"01",x"39",x"81",x"BA",x"27",
    x"A4",x"81",x"2C",x"27",x"54",x"81",x"3B",x"27",x"5F",x"81",x"BE",x"27",x"68",x"8D",x"79",x"34",
    x"02",x"BD",x"D6",x"C4",x"27",x"0E",x"B6",x"2C",x"36",x"27",x"09",x"9B",x"51",x"B1",x"2C",x"37",
    x"23",x"02",x"8D",x"29",x"8D",x"7E",x"35",x"02",x"8D",x"6C",x"27",x"06",x"8D",x"1F",x"9D",x"C6",
    x"20",x"C8",x"4D",x"27",x"08",x"9D",x"C6",x"81",x"2C",x"27",x"02",x"8D",x"7A",x"9D",x"C6",x"26",
    x"BC",x"20",x"0A",x"BD",x"D6",x"C4",x"27",x"05",x"B6",x"2C",x"36",x"27",x"AF",x"86",x"0D",x"8D",
    x"68",x"8D",x"43",x"26",x"A7",x"86",x"0A",x"20",x"60",x"BD",x"D6",x"C4",x"27",x"0C",x"F6",x"2C",
    x"36",x"F1",x"2C",x"35",x"25",x"07",x"8D",x"E5",x"20",x"1A",x"F6",x"2C",x"36",x"F0",x"2C",x"34",
    x"24",x"FB",x"50",x"20",x"09",x"BD",x"C1",x"4C",x"81",x"29",x"10",x"26",x"F5",x"E6",x"8D",x"16",
    x"26",x"02",x"8D",x"1C",x"9D",x"C0",x"20",x"A8",x"BD",x"B9",x"06",x"BD",x"B9",x"45",x"27",x"05",
    x"BD",x"BF",x"89",x"86",x"FF",x"39",x"BD",x"D6",x"C4",x"7D",x"29",x"4D",x"39",x"8D",x"18",x"5A",
    x"5D",x"26",x"FA",x"39",x"D6",x"51",x"8E",x"23",x"2F",x"5C",x"5A",x"27",x"15",x"A6",x"80",x"8D",
    x"08",x"20",x"F7",x"86",x"3F",x"8D",x"02",x"86",x"20",x"7E",x"D6",x"A2",x"8D",x"FB",x"A6",x"80",
    x"26",x"FA",x"39",x"35",x"10",x"8D",x"F7",x"6E",x"84",x"27",x"82",x"8D",x"03",x"0F",x"77",x"39",
    x"81",x"23",x"26",x"07",x"BD",x"C2",x"72",x"27",x"F0",x"9D",x"BA",x"8D",x"AB",x"27",x"12",x"8D",
    x"C3",x"9D",x"C6",x"27",x"E4",x"86",x"2C",x"8D",x"AD",x"27",x"02",x"86",x"0D",x"8D",x"10",x"20",
    x"E8",x"8D",x"06",x"8D",x"AF",x"8D",x"02",x"20",x"E8",x"8D",x"9B",x"26",x"D2",x"86",x"22",x"20",
    x"B8",x"BD",x"B8",x"DA",x"BD",x"B9",x"06",x"C6",x"01",x"34",x"04",x"BD",x"B9",x"45",x"27",x"0C",
    x"BD",x"C1",x"55",x"E7",x"E4",x"10",x"27",x"FB",x"9A",x"BD",x"BF",x"2E",x"35",x"04",x"D7",x"66",
    x"BD",x"BF",x"4A",x"D6",x"66",x"34",x"04",x"9D",x"BA",x"BD",x"B8",x"D5",x"35",x"04",x"D7",x"66",
    x"20",x"14",x"30",x"E4",x"D6",x"66",x"3A",x"BD",x"BE",x"75",x"5C",x"5A",x"27",x"15",x"A6",x"80",
    x"A1",x"C0",x"27",x"F7",x"0C",x"66",x"E6",x"E4",x"D0",x"66",x"25",x"05",x"5C",x"D1",x"51",x"24",
    x"E1",x"0F",x"66",x"BD",x"BE",x"CB",x"D6",x"66",x"7E",x"BD",x"D6",x"9D",x"C0",x"BD",x"B8",x"DA",
    x"BD",x"BB",x"7C",x"34",x"12",x"E6",x"84",x"34",x"04",x"BD",x"DC",x"23",x"BD",x"C1",x"60",x"D7",
    x"6A",x"10",x"27",x"FB",x"3E",x"C6",x"FF",x"81",x"29",x"27",x"03",x"BD",x"C1",x"60",x"D7",x"69",
    x"BD",x"B8",x"D7",x"C6",x"D4",x"9D",x"BD",x"BD",x"BF",x"30",x"A6",x"E0",x"90",x"6A",x"10",x"25",
    x"FB",x"21",x"4C",x"91",x"69",x"24",x"02",x"97",x"69",x"96",x"69",x"26",x"02",x"35",x"92",x"91",
    x"51",x"24",x"04",x"96",x"69",x"97",x"51",x"35",x"12",x"BD",x"DC",x"27",x"AE",x"01",x"D6",x"6A",
    x"5A",x"3A",x"BD",x"BE",x"37",x"7E",x"DC",x"23",x"DD",x"50",x"BD",x"B8",x"8B",x"BD",x"BF",x"7F",
    x"30",x"01",x"39",x"8E",x"C4",x"CA",x"8D",x"04",x"DC",x"31",x"8D",x"EC",x"7E",x"C3",x"4E",x"0D",
    x"77",x"26",x"EF",x"7E",x"D9",x"A3",x"BD",x"C2",x"DD",x"BD",x"D9",x"2F",x"96",x"6D",x"9C",x"6E",
    x"26",x"0F",x"90",x"70",x"26",x"0B",x"F6",x"2C",x"44",x"32",x"EB",x"BD",x"D3",x"4F",x"7E",x"B6",
    x"AB",x"9F",x"6B",x"EC",x"84",x"27",x"37",x"BD",x"CE",x"EC",x"BD",x"CC",x"BB",x"26",x"27",x"9E",
    x"6B",x"EC",x"02",x"FD",x"2C",x"40",x"8D",x"C2",x"8E",x"29",x"5B",x"86",x"20",x"BD",x"D6",x"A2",
    x"A6",x"80",x"27",x"0D",x"2A",x"F7",x"BD",x"E8",x"1A",x"BD",x"C3",x"47",x"BD",x"E8",x"1A",x"20",
    x"EF",x"8D",x"AC",x"BD",x"C2",x"DD",x"9E",x"6B",x"EC",x"84",x"30",x"8B",x"20",x"AB",x"8E",x"60",
    x"01",x"0C",x"6D",x"96",x"6D",x"BD",x"DC",x"19",x"20",x"9F",x"20",x"49",x"6E",x"20",x"00",x"4F",
    x"5F",x"DD",x"6B",x"43",x"53",x"FD",x"2C",x"3C",x"8E",x"F9",x"FF",x"9F",x"6E",x"8D",x"63",x"27",
    x"1C",x"8D",x"4F",x"9F",x"6B",x"8D",x"5B",x"26",x"04",x"9F",x"6E",x"20",x"10",x"C6",x"C8",x"9D",
    x"BD",x"8D",x"4F",x"27",x"08",x"8D",x"3B",x"8D",x"49",x"26",x"34",x"9F",x"6E",x"81",x"2C",x"26",
    x"07",x"9D",x"C0",x"8D",x"38",x"BF",x"2C",x"3C",x"9E",x"6E",x"34",x"10",x"9C",x"6B",x"25",x"42",
    x"30",x"01",x"9F",x"33",x"BD",x"B3",x"E6",x"9F",x"6E",x"97",x"70",x"9E",x"6B",x"34",x"10",x"9F",
    x"33",x"BD",x"B3",x"E6",x"9F",x"6B",x"97",x"6D",x"35",x"60",x"39",x"9D",x"C6",x"27",x"FB",x"7E",
    x"B8",x"F4",x"81",x"2E",x"26",x"07",x"BE",x"2C",x"40",x"9F",x"33",x"0E",x"C0",x"BD",x"CA",x"25",
    x"0E",x"C6",x"9D",x"C6",x"27",x"02",x"81",x"2C",x"39",x"81",x"41",x"25",x"04",x"80",x"5B",x"80",
    x"A5",x"39",x"7E",x"BF",x"43",x"C6",x"03",x"8C",x"C6",x"02",x"8C",x"C6",x"04",x"8C",x"C6",x"08",
    x"34",x"04",x"BD",x"C5",x"49",x"25",x"C8",x"34",x"02",x"1F",x"89",x"9D",x"C0",x"81",x"C8",x"26",
    x"0B",x"9D",x"C0",x"1F",x"89",x"BD",x"C5",x"49",x"25",x"B5",x"9D",x"C0",x"1F",x"98",x"E6",x"E4",
    x"A0",x"E0",x"25",x"AB",x"8E",x"2B",x"29",x"3A",x"35",x"04",x"E7",x"80",x"4A",x"2A",x"FB",x"9D",
    x"C6",x"27",x"97",x"34",x"04",x"9D",x"BA",x"20",x"C9",x"27",x"B7",x"8D",x"03",x"7E",x"B6",x"AB",
    x"8D",x"A0",x"34",x"01",x"BD",x"C4",x"CF",x"35",x"01",x"26",x"01",x"39",x"BD",x"D2",x"03",x"9E",
    x"6B",x"DE",x"6E",x"96",x"70",x"BD",x"DC",x"19",x"4F",x"5F",x"1F",x"12",x"33",x"CB",x"EC",x"C4",
    x"27",x"18",x"30",x"AB",x"8C",x"9F",x"FC",x"25",x"F1",x"BD",x"DC",x"2D",x"BD",x"D5",x"F3",x"63",
    x"84",x"8E",x"60",x"01",x"9F",x"6B",x"0C",x"6D",x"20",x"D2",x"BD",x"DC",x"2D",x"BD",x"D5",x"F3",
    x"96",x"70",x"91",x"21",x"27",x"0B",x"63",x"84",x"0C",x"70",x"8E",x"60",x"01",x"9F",x"6E",x"20",
    x"BB",x"96",x"6D",x"7E",x"B3",x"B9",x"54",x"52",x"41",x"BD",x"D2",x"09",x"8D",x"2A",x"03",x"72",
    x"9D",x"C6",x"81",x"22",x"26",x"17",x"CE",x"C5",x"F6",x"BD",x"D1",x"AD",x"0C",x"77",x"73",x"22",
    x"4D",x"73",x"28",x"17",x"7C",x"22",x"4C",x"BD",x"D4",x"1D",x"BD",x"B8",x"E7",x"BD",x"C4",x"CF",
    x"10",x"BF",x"2C",x"38",x"FF",x"2C",x"3A",x"39",x"0F",x"72",x"C6",x"12",x"7E",x"D3",x"51",x"BD",
    x"D2",x"09",x"8E",x"00",x"0A",x"81",x"2C",x"27",x"07",x"9D",x"C6",x"27",x"03",x"BD",x"CA",x"25",
    x"BF",x"2C",x"46",x"8E",x"00",x"0A",x"9D",x"C6",x"27",x"0E",x"9D",x"BA",x"27",x"0D",x"BD",x"CA",
    x"25",x"10",x"27",x"F8",x"EE",x"BD",x"C5",x"2B",x"BF",x"2C",x"48",x"7C",x"2C",x"45",x"32",x"62",
    x"7E",x"B2",x"A8",x"F6",x"2C",x"45",x"27",x"BF",x"BE",x"2C",x"46",x"BD",x"CB",x"9E",x"25",x"17",
    x"73",x"2C",x"45",x"BD",x"C3",x"53",x"4C",x"69",x"6E",x"65",x"20",x"6E",x"6F",x"74",x"20",x"65",
    x"6D",x"70",x"74",x"79",x"0D",x"0A",x"00",x"FC",x"2C",x"46",x"BD",x"C4",x"48",x"34",x"10",x"A6",
    x"80",x"26",x"FC",x"86",x"20",x"A7",x"1F",x"6F",x"84",x"35",x"10",x"BD",x"E0",x"79",x"25",x"25",
    x"9F",x"C7",x"9D",x"C0",x"24",x"1F",x"BD",x"CA",x"25",x"1F",x"10",x"F3",x"2C",x"48",x"FD",x"2C",
    x"46",x"C6",x"06",x"10",x"25",x"5B",x"00",x"B6",x"2C",x"45",x"2A",x"0C",x"73",x"2C",x"45",x"9D",
    x"C6",x"27",x"A0",x"20",x"03",x"7F",x"2C",x"45",x"8E",x"29",x"5A",x"32",x"62",x"7E",x"B2",x"B0",
    x"86",x"01",x"97",x"7B",x"34",x"02",x"5A",x"BD",x"C8",x"83",x"9D",x"C6",x"26",x"05",x"35",x"02",
    x"7E",x"C7",x"73",x"D7",x"80",x"BD",x"BF",x"30",x"D1",x"7B",x"23",x"04",x"D6",x"7B",x"D7",x"51",
    x"BD",x"C3",x"34",x"35",x"02",x"81",x"26",x"27",x"07",x"D6",x"7B",x"D0",x"51",x"BD",x"C3",x"30",
    x"7E",x"C8",x"61",x"D7",x"80",x"9F",x"0A",x"86",x"02",x"97",x"7B",x"A6",x"84",x"81",x"25",x"27",
    x"C3",x"81",x"20",x"26",x"07",x"0C",x"7B",x"30",x"01",x"5A",x"26",x"EF",x"9E",x"0A",x"D6",x"80",
    x"86",x"25",x"BD",x"C8",x"83",x"BD",x"D6",x"A2",x"20",x"21",x"9D",x"C0",x"BD",x"BF",x"30",x"BD",
    x"BF",x"4A",x"C6",x"3B",x"9D",x"BD",x"30",x"E4",x"9F",x"7D",x"20",x"06",x"96",x"7F",x"27",x"08",
    x"9E",x"7D",x"0F",x"7F",x"E6",x"80",x"26",x"03",x"7E",x"BF",x"43",x"0F",x"7C",x"0F",x"7B",x"A6",
    x"80",x"81",x"21",x"10",x"27",x"FF",x"79",x"81",x"26",x"26",x"05",x"03",x"7B",x"7E",x"C6",x"D4",
    x"81",x"23",x"27",x"65",x"5A",x"26",x"15",x"BD",x"C8",x"83",x"BD",x"D6",x"A2",x"9D",x"C6",x"26",
    x"CB",x"96",x"7F",x"26",x"03",x"BD",x"C2",x"D3",x"BD",x"BE",x"C7",x"39",x"81",x"2B",x"26",x"09",
    x"BD",x"C8",x"83",x"86",x"08",x"97",x"7C",x"20",x"C4",x"81",x"2E",x"27",x"59",x"81",x"25",x"10",
    x"27",x"FF",x"70",x"81",x"3D",x"26",x"07",x"A6",x"80",x"5A",x"27",x"CB",x"20",x"84",x"A1",x"84",
    x"26",x"FA",x"81",x"24",x"27",x"19",x"81",x"2A",x"26",x"F2",x"96",x"7C",x"8A",x"20",x"97",x"7C",
    x"C1",x"02",x"25",x"11",x"A6",x"01",x"81",x"24",x"26",x"0B",x"5A",x"30",x"01",x"0C",x"7B",x"96",
    x"7C",x"8A",x"10",x"97",x"7C",x"30",x"01",x"0C",x"7B",x"0F",x"7A",x"0C",x"7B",x"5A",x"27",x"47",
    x"A6",x"80",x"81",x"2E",x"27",x"1C",x"81",x"23",x"27",x"F1",x"81",x"2C",x"26",x"1F",x"96",x"7C",
    x"8A",x"40",x"97",x"7C",x"20",x"E5",x"A6",x"84",x"81",x"23",x"26",x"B0",x"86",x"01",x"97",x"7A",
    x"30",x"01",x"0C",x"7A",x"5A",x"27",x"20",x"A6",x"80",x"81",x"23",x"27",x"F5",x"81",x"5E",x"26",
    x"16",x"A1",x"84",x"26",x"12",x"A1",x"01",x"26",x"0E",x"A1",x"02",x"26",x"0A",x"C1",x"04",x"25",
    x"06",x"C0",x"04",x"30",x"04",x"0C",x"7C",x"30",x"1F",x"0C",x"7B",x"96",x"7C",x"85",x"08",x"26",
    x"18",x"0A",x"7B",x"5D",x"27",x"13",x"A6",x"84",x"80",x"2D",x"27",x"06",x"81",x"FE",x"26",x"09",
    x"86",x"08",x"8A",x"04",x"9A",x"7C",x"97",x"7C",x"5A",x"9D",x"C6",x"10",x"27",x"FF",x"34",x"D7",
    x"80",x"BD",x"B8",x"F8",x"96",x"7B",x"9B",x"7A",x"81",x"19",x"10",x"24",x"FE",x"FA",x"96",x"7C",
    x"8A",x"80",x"97",x"7C",x"10",x"8E",x"2B",x"A7",x"CE",x"C5",x"18",x"BD",x"B0",x"02",x"BD",x"C3",
    x"4E",x"0F",x"7F",x"9D",x"C6",x"27",x"0C",x"97",x"7F",x"81",x"3B",x"27",x"04",x"9D",x"BA",x"20",
    x"02",x"9D",x"C0",x"9E",x"7D",x"E6",x"80",x"D0",x"80",x"3A",x"D6",x"80",x"10",x"26",x"FE",x"CB",
    x"7E",x"C7",x"6D",x"34",x"02",x"86",x"2B",x"0D",x"7C",x"27",x"03",x"BD",x"D6",x"A2",x"35",x"82",
    x"9D",x"C0",x"C6",x"87",x"9D",x"BD",x"C6",x"BB",x"9D",x"BD",x"BD",x"CA",x"25",x"27",x"11",x"BD",
    x"B3",x"E6",x"10",x"25",x"EE",x"2C",x"B7",x"2C",x"31",x"BF",x"2C",x"2F",x"7E",x"DC",x"23",x"39",
    x"BF",x"2C",x"2F",x"B6",x"2C",x"29",x"27",x"F7",x"BE",x"2C",x"2A",x"9F",x"31",x"7E",x"B2",x"36",
    x"BD",x"C1",x"4E",x"26",x"EA",x"5D",x"26",x"0A",x"7E",x"BF",x"43",x"F6",x"2C",x"29",x"26",x"04",
    x"C6",x"14",x"0E",x"B7",x"5F",x"F7",x"2C",x"26",x"81",x"82",x"27",x"27",x"9D",x"C6",x"24",x"0A",
    x"BD",x"B7",x"8E",x"26",x"1D",x"BD",x"B6",x"8D",x"20",x"15",x"BD",x"C5",x"2D",x"FE",x"2C",x"2A",
    x"BE",x"2C",x"2C",x"B6",x"2C",x"2E",x"DF",x"31",x"9F",x"C7",x"97",x"1A",x"BD",x"DC",x"19",x"7F",
    x"2C",x"29",x"39",x"9D",x"C0",x"8D",x"E3",x"6D",x"80",x"26",x"02",x"30",x"03",x"9F",x"C7",x"7E",
    x"B6",x"E4",x"BD",x"B8",x"DA",x"BD",x"BB",x"96",x"9F",x"50",x"BD",x"DC",x"14",x"BD",x"C1",x"F9",
    x"BD",x"BD",x"D9",x"BD",x"DC",x"23",x"7E",x"B8",x"D7",x"81",x"FF",x"10",x"27",x"11",x"BA",x"81",
    x"BD",x"10",x"27",x"23",x"CE",x"81",x"C0",x"10",x"26",x"5E",x"67",x"8D",x"0C",x"34",x"10",x"C6",
    x"D4",x"9D",x"BD",x"BD",x"C1",x"66",x"AF",x"F1",x"39",x"5F",x"9D",x"C0",x"24",x"06",x"80",x"30",
    x"1F",x"89",x"9D",x"C0",x"8E",x"27",x"AA",x"58",x"3A",x"39",x"8D",x"ED",x"34",x"10",x"BD",x"B8",
    x"D3",x"BD",x"C1",x"E1",x"8E",x"21",x"4E",x"BD",x"B9",x"45",x"26",x"07",x"BD",x"BE",x"75",x"E7",
    x"84",x"EF",x"01",x"96",x"05",x"EE",x"F1",x"BD",x"B0",x"0E",x"97",x"05",x"BD",x"B9",x"45",x"26",
    x"0C",x"E6",x"84",x"D7",x"51",x"AE",x"01",x"CE",x"23",x"2F",x"BD",x"DC",x"01",x"7E",x"DC",x"23",
    x"80",x"C3",x"27",x"0B",x"81",x"D3",x"26",x"0C",x"7D",x"2B",x"37",x"27",x"07",x"8D",x"08",x"B7",
    x"2B",x"3B",x"0E",x"C0",x"7E",x"B8",x"F4",x"34",x"01",x"1A",x"50",x"BE",x"2B",x"35",x"BF",x"23",
    x"0F",x"7F",x"2B",x"34",x"35",x"81",x"9D",x"C0",x"C6",x"D4",x"9D",x"BD",x"BD",x"BA",x"A2",x"BF",
    x"2B",x"35",x"10",x"27",x"F5",x"7D",x"C6",x"FF",x"8E",x"2B",x"37",x"20",x"25",x"9D",x"C0",x"C6",
    x"D4",x"9D",x"BD",x"BD",x"E3",x"EB",x"86",x"0A",x"8E",x"2B",x"69",x"30",x"1C",x"E1",x"84",x"27",
    x"11",x"4A",x"26",x"F7",x"86",x"0A",x"6D",x"84",x"27",x"08",x"30",x"04",x"4A",x"26",x"F7",x"7E",
    x"B1",x"FC",x"E7",x"84",x"C6",x"87",x"9D",x"BD",x"80",x"BB",x"27",x"08",x"81",x"01",x"10",x"26",
    x"EE",x"F2",x"86",x"80",x"34",x"12",x"9D",x"C0",x"8D",x"1B",x"27",x"14",x"BD",x"B3",x"E6",x"10",
    x"25",x"EC",x"BF",x"AA",x"E0",x"35",x"40",x"30",x"1F",x"AF",x"41",x"A7",x"43",x"7E",x"DC",x"23",
    x"35",x"42",x"6F",x"C4",x"39",x"9D",x"C6",x"BD",x"B7",x"8E",x"9E",x"33",x"39",x"7E",x"BF",x"43",
    x"BD",x"D2",x"09",x"BD",x"B4",x"3F",x"CC",x"00",x"0A",x"DD",x"D8",x"DD",x"DA",x"5F",x"DD",x"DC",
    x"4A",x"DD",x"DE",x"9D",x"C6",x"24",x"04",x"8D",x"DC",x"9F",x"D8",x"BD",x"B8",x"E7",x"27",x"04",
    x"8D",x"D3",x"9F",x"DC",x"BD",x"B8",x"E7",x"27",x"08",x"8D",x"CA",x"9C",x"DC",x"25",x"CE",x"9F",
    x"DE",x"BD",x"B8",x"E7",x"27",x"06",x"8D",x"BD",x"9F",x"DA",x"27",x"C1",x"BD",x"C5",x"2B",x"8D",
    x"16",x"BD",x"CB",x"A3",x"8D",x"10",x"BD",x"B4",x"3F",x"7E",x"B2",x"9B",x"A6",x"80",x"A7",x"A0",
    x"81",x"20",x"27",x"F8",x"0E",x"CD",x"86",x"4F",x"97",x"E2",x"BD",x"B4",x"20",x"30",x"01",x"BD",
    x"CF",x"EC",x"26",x"01",x"39",x"DF",x"31",x"30",x"1D",x"9F",x"E0",x"30",x"04",x"10",x"8E",x"29",
    x"58",x"EF",x"A1",x"0F",x"E3",x"8D",x"D5",x"4D",x"27",x"17",x"2A",x"F9",x"C6",x"0D",x"CE",x"CC",
    x"7C",x"A1",x"C5",x"27",x"05",x"5A",x"2A",x"F9",x"20",x"EB",x"58",x"CB",x"0E",x"AD",x"D5",x"20",
    x"E6",x"0D",x"E3",x"27",x"07",x"1F",x"20",x"83",x"29",x"56",x"8D",x"08",x"9E",x"E0",x"EC",x"84",
    x"30",x"8B",x"20",x"BB",x"34",x"06",x"96",x"1A",x"9E",x"E0",x"7E",x"B3",x"01",x"8D",x"9D",x"81",
    x"87",x"26",x"18",x"86",x"4F",x"97",x"4E",x"8D",x"93",x"81",x"BB",x"27",x"04",x"81",x"BC",x"26",
    x"0A",x"8D",x"09",x"81",x"2C",x"27",x"FA",x"81",x"C8",x"27",x"F6",x"39",x"BD",x"CA",x"7C",x"30",
    x"1F",x"31",x"3F",x"9F",x"C7",x"24",x"40",x"34",x"30",x"BD",x"B7",x"8E",x"8D",x"5E",x"25",x"20",
    x"0D",x"E2",x"27",x"1C",x"EC",x"C4",x"26",x"04",x"96",x"4E",x"26",x"14",x"EC",x"42",x"81",x"FF",
    x"27",x"28",x"DD",x"50",x"BD",x"B8",x"8B",x"BD",x"BF",x"7F",x"0C",x"E3",x"30",x"01",x"AF",x"E4",
    x"35",x"30",x"BD",x"CA",x"7C",x"25",x"FB",x"9E",x"C7",x"31",x"3F",x"A6",x"82",x"81",x"20",x"26",
    x"04",x"A7",x"A0",x"20",x"F6",x"9E",x"C7",x"7E",x"CA",x"7C",x"34",x"40",x"BD",x"C3",x"53",x"55",
    x"6E",x"64",x"65",x"66",x"69",x"6E",x"65",x"64",x"20",x"4C",x"69",x"6E",x"65",x"20",x"00",x"EC",
    x"F1",x"BD",x"C4",x"5A",x"BD",x"C4",x"53",x"BD",x"C2",x"DD",x"20",x"C4",x"DC",x"33",x"10",x"93",
    x"DC",x"25",x"27",x"10",x"93",x"DE",x"22",x"22",x"DE",x"1B",x"20",x"07",x"10",x"A3",x"C4",x"27",
    x"1B",x"33",x"44",x"11",x"93",x"1D",x"26",x"F4",x"0D",x"E2",x"26",x"0E",x"ED",x"C1",x"CC",x"FF",
    x"FF",x"ED",x"C1",x"DF",x"1D",x"1F",x"30",x"BD",x"B1",x"E5",x"43",x"39",x"4F",x"39",x"9F",x"33",
    x"7E",x"B3",x"E6",x"9E",x"DC",x"8D",x"F7",x"34",x"12",x"9E",x"D8",x"8D",x"F1",x"A1",x"E4",x"22",
    x"06",x"25",x"68",x"AC",x"61",x"25",x"64",x"32",x"63",x"8D",x"01",x"86",x"4F",x"97",x"E2",x"DC",
    x"D8",x"DD",x"50",x"9E",x"DC",x"8D",x"D7",x"97",x"1A",x"EC",x"84",x"26",x"10",x"A6",x"02",x"27",
    x"19",x"0C",x"1A",x"96",x"1A",x"BD",x"DC",x"19",x"8E",x"60",x"01",x"20",x"EC",x"EC",x"02",x"10",
    x"93",x"DE",x"23",x"07",x"D3",x"DA",x"93",x"50",x"23",x"31",x"39",x"0D",x"E2",x"27",x"1B",x"10",
    x"9E",x"50",x"10",x"AF",x"02",x"DE",x"1B",x"20",x"07",x"10",x"A3",x"C4",x"27",x"09",x"33",x"44",
    x"11",x"93",x"1D",x"26",x"F4",x"20",x"03",x"10",x"AF",x"42",x"EC",x"84",x"30",x"8B",x"DC",x"50",
    x"D3",x"DA",x"DD",x"50",x"25",x"05",x"83",x"FA",x"00",x"25",x"AE",x"7E",x"BF",x"43",x"C6",x"FF",
    x"5C",x"BD",x"CA",x"7C",x"81",x"D4",x"27",x"F8",x"81",x"D5",x"27",x"F4",x"81",x"D3",x"27",x"F0",
    x"30",x"1F",x"31",x"3F",x"5D",x"10",x"26",x"FE",x"C3",x"39",x"BD",x"CA",x"7C",x"27",x"FA",x"81",
    x"87",x"26",x"F7",x"7E",x"CA",x"E3",x"BD",x"CA",x"7C",x"30",x"1F",x"31",x"3F",x"81",x"22",x"10",
    x"26",x"FE",x"9E",x"5F",x"BD",x"CA",x"7C",x"10",x"27",x"FE",x"98",x"81",x"2C",x"26",x"03",x"5D",
    x"27",x"F5",x"81",x"22",x"26",x"0A",x"BD",x"CA",x"7C",x"4D",x"27",x"EB",x"81",x"22",x"26",x"F6",
    x"81",x"28",x"26",x"01",x"5C",x"81",x"29",x"26",x"01",x"5A",x"20",x"D8",x"8A",x"99",x"C4",x"8F",
    x"88",x"FF",x"87",x"98",x"C1",x"B0",x"F4",x"AD",x"9B",x"F6",x"CA",x"FC",x"CA",x"FC",x"CA",x"FC",
    x"CA",x"FC",x"CA",x"FC",x"CA",x"7C",x"CA",x"E4",x"CA",x"DD",x"CC",x"1E",x"CC",x"3A",x"CC",x"53",
    x"CC",x"46",x"CA",x"F1",x"CC",x"53",x"BD",x"BF",x"30",x"BD",x"BF",x"4A",x"35",x"04",x"10",x"FF",
    x"2C",x"42",x"F7",x"2C",x"44",x"BD",x"B8",x"E7",x"7E",x"D1",x"C6",x"34",x"76",x"8E",x"29",x"5A",
    x"F6",x"2C",x"44",x"27",x"12",x"FE",x"2C",x"42",x"30",x"01",x"31",x"84",x"A6",x"A0",x"27",x"09",
    x"A1",x"C0",x"26",x"EC",x"5A",x"26",x"F5",x"35",x"F6",x"43",x"35",x"F6",x"9D",x"C0",x"C6",x"A1",
    x"9D",x"BD",x"8D",x"28",x"17",x"00",x"7E",x"0F",x"77",x"BD",x"BB",x"96",x"9F",x"48",x"97",x"4A",
    x"BD",x"BF",x"38",x"8E",x"29",x"5A",x"4F",x"BD",x"BF",x"92",x"7E",x"B7",x"D8",x"9D",x"C0",x"D6",
    x"08",x"26",x"07",x"F6",x"2B",x"D6",x"10",x"26",x"F6",x"39",x"39",x"C6",x"5F",x"F7",x"2B",x"D6",
    x"0F",x"08",x"BD",x"C1",x"22",x"81",x"3B",x"26",x"02",x"9D",x"C0",x"81",x"23",x"26",x"0A",x"BD",
    x"D3",x"A7",x"BD",x"D6",x"FC",x"03",x"08",x"9D",x"BA",x"81",x"22",x"26",x"D2",x"BD",x"B8",x"5B",
    x"0D",x"08",x"26",x"03",x"BD",x"C3",x"34",x"9D",x"C6",x"81",x"3B",x"27",x"C0",x"0E",x"BA",x"9E",
    x"3C",x"9F",x"31",x"7E",x"B8",x"F4",x"9F",x"C7",x"BD",x"B6",x"EC",x"6D",x"80",x"26",x"0B",x"C6",
    x"04",x"BD",x"CF",x"EC",x"27",x"28",x"DF",x"3C",x"30",x"01",x"9F",x"C7",x"9D",x"C6",x"81",x"83",
    x"26",x"E6",x"7E",x"CE",x"4B",x"BD",x"E0",x"76",x"CC",x"00",x"00",x"FD",x"23",x"20",x"B6",x"22",
    x"A9",x"F7",x"22",x"A9",x"10",x"25",x"E7",x"A9",x"0D",x"78",x"27",x"8E",x"C6",x"36",x"0E",x"B7",
    x"9D",x"C0",x"81",x"B8",x"10",x"27",x"0D",x"16",x"81",x"F3",x"10",x"27",x"0D",x"03",x"81",x"F8",
    x"10",x"27",x"21",x"B0",x"81",x"97",x"26",x"25",x"9D",x"C0",x"BD",x"CA",x"25",x"BF",x"29",x"54",
    x"C6",x"3B",x"9D",x"BD",x"BD",x"C1",x"4E",x"86",x"32",x"3D",x"FD",x"23",x"20",x"10",x"27",x"F1",
    x"92",x"9D",x"BA",x"F7",x"2B",x"D6",x"0F",x"08",x"BD",x"CD",x"29",x"20",x"03",x"BD",x"CD",x"0B",
    x"4F",x"BD",x"D6",x"F1",x"2B",x"0E",x"8D",x"9D",x"BE",x"29",x"54",x"9F",x"33",x"4D",x"10",x"26",
    x"E8",x"BB",x"86",x"2C",x"8E",x"29",x"5A",x"A7",x"84",x"5F",x"20",x"33",x"C6",x"3A",x"BD",x"D6",
    x"F1",x"26",x"9B",x"96",x"08",x"10",x"26",x"FF",x"56",x"BD",x"C3",x"53",x"3F",x"52",x"65",x"64",
    x"6F",x"20",x"66",x"72",x"6F",x"6D",x"20",x"73",x"74",x"61",x"72",x"74",x"0D",x"0A",x"00",x"9E",
    x"38",x"9F",x"C7",x"96",x"35",x"97",x"1A",x"7E",x"DC",x"19",x"9E",x"3E",x"D6",x"40",x"86",x"4F",
    x"97",x"08",x"9F",x"41",x"D7",x"43",x"8C",x"9D",x"BA",x"BD",x"BB",x"96",x"9F",x"48",x"97",x"4A",
    x"9E",x"C7",x"96",x"1A",x"9F",x"33",x"97",x"35",x"9E",x"41",x"96",x"43",x"8D",x"D7",x"A6",x"84",
    x"9D",x"CD",x"26",x"15",x"96",x"08",x"10",x"26",x"FF",x"0C",x"BD",x"D6",x"F1",x"27",x"9D",x"2A",
    x"05",x"BD",x"EB",x"3B",x"20",x"03",x"BD",x"CD",x"65",x"9F",x"C7",x"BD",x"B9",x"45",x"27",x"67",
    x"9D",x"C0",x"10",x"9E",x"C7",x"96",x"05",x"34",x"22",x"CE",x"C4",x"0A",x"81",x"08",x"26",x"04",
    x"33",x"C9",x"FF",x"FB",x"BD",x"B0",x"02",x"35",x"02",x"10",x"AC",x"E1",x"27",x"CF",x"10",x"9F",
    x"C7",x"BD",x"B0",x"27",x"CE",x"B0",x"2C",x"96",x"8B",x"34",x"02",x"AD",x"C4",x"35",x"02",x"BD",
    x"DC",x"27",x"9D",x"C6",x"27",x"06",x"81",x"2C",x"10",x"26",x"FF",x"50",x"9E",x"C7",x"9F",x"41",
    x"96",x"1A",x"97",x"43",x"9E",x"33",x"9F",x"C7",x"BD",x"CE",x"03",x"9D",x"C6",x"10",x"26",x"FF",
    x"76",x"9E",x"41",x"D6",x"08",x"27",x"07",x"96",x"43",x"97",x"40",x"9F",x"3E",x"39",x"A6",x"84",
    x"10",x"26",x"FF",x"35",x"0F",x"77",x"39",x"4F",x"5F",x"BD",x"D6",x"C4",x"7D",x"29",x"4D",x"26",
    x"1E",x"9D",x"C0",x"9E",x"C7",x"1F",x"89",x"81",x"22",x"27",x"14",x"30",x"1F",x"CC",x"3A",x"2C",
    x"8D",x"14",x"0C",x"51",x"0A",x"51",x"27",x"06",x"A6",x"82",x"81",x"20",x"27",x"F6",x"8C",x"8D",
    x"05",x"CE",x"B7",x"D8",x"20",x"91",x"BD",x"BF",x"94",x"9F",x"C7",x"39",x"BD",x"27",x"DC",x"BD",
    x"D2",x"09",x"CE",x"D4",x"2A",x"7E",x"B0",x"02",x"30",x"01",x"8C",x"9E",x"C7",x"8D",x"06",x"8E",
    x"29",x"59",x"9F",x"C7",x"39",x"BD",x"27",x"D6",x"CE",x"29",x"5A",x"0F",x"DA",x"0F",x"DB",x"A6",
    x"80",x"27",x"21",x"0D",x"DA",x"27",x"0F",x"BD",x"CF",x"D1",x"24",x"18",x"81",x"30",x"25",x"04",
    x"81",x"39",x"23",x"10",x"0F",x"DA",x"81",x"20",x"27",x"0A",x"97",x"D9",x"81",x"22",x"27",x"35",
    x"0D",x"DB",x"27",x"16",x"A7",x"C0",x"27",x"06",x"81",x"3A",x"27",x"CF",x"20",x"D1",x"6F",x"C0",
    x"6F",x"C0",x"6F",x"C4",x"1F",x"30",x"83",x"29",x"58",x"39",x"81",x"3F",x"26",x"04",x"86",x"AB",
    x"20",x"E2",x"81",x"27",x"26",x"13",x"CC",x"3A",x"8D",x"ED",x"C1",x"0F",x"D9",x"A6",x"80",x"27",
    x"D3",x"91",x"D9",x"27",x"CF",x"A7",x"C0",x"20",x"F4",x"81",x"30",x"25",x"04",x"81",x"3C",x"25",
    x"C3",x"30",x"1F",x"34",x"40",x"0F",x"D8",x"CE",x"27",x"66",x"5F",x"D7",x"D9",x"33",x"4A",x"E6",
    x"C4",x"27",x"37",x"10",x"AE",x"41",x"34",x"40",x"CE",x"D4",x"97",x"BD",x"B0",x"02",x"35",x"40",
    x"E1",x"C4",x"25",x"04",x"DB",x"D9",x"20",x"E3",x"DB",x"D9",x"CA",x"80",x"35",x"40",x"96",x"D8",
    x"26",x"06",x"C1",x"8F",x"26",x"06",x"86",x"3A",x"ED",x"C1",x"20",x"90",x"E7",x"C0",x"C1",x"83",
    x"26",x"02",x"0C",x"DB",x"C1",x"8C",x"27",x"A3",x"20",x"F0",x"CE",x"27",x"6B",x"03",x"D8",x"26",
    x"B9",x"35",x"40",x"A6",x"80",x"A7",x"C0",x"8D",x"08",x"25",x"DF",x"03",x"DA",x"A7",x"5F",x"20",
    x"D9",x"81",x"61",x"25",x"06",x"81",x"7A",x"22",x"02",x"88",x"20",x"7E",x"C5",x"49",x"D8",x"C4",
    x"C1",x"F5",x"EE",x"91",x"EE",x"8A",x"EE",x"A9",x"EE",x"59",x"EE",x"98",x"EE",x"81",x"26",x"10",
    x"A6",x"84",x"27",x"10",x"0C",x"1A",x"96",x"1A",x"BD",x"DC",x"19",x"8E",x"60",x"01",x"20",x"EC",
    x"EE",x"80",x"9F",x"C7",x"39",x"10",x"DF",x"75",x"BD",x"D9",x"0A",x"9E",x"C7",x"9F",x"38",x"A6",
    x"80",x"27",x"07",x"81",x"3A",x"27",x"2E",x"7E",x"B8",x"F4",x"8D",x"D0",x"27",x"72",x"DF",x"31",
    x"96",x"72",x"27",x"21",x"11",x"B3",x"2C",x"38",x"25",x"1B",x"11",x"B3",x"2C",x"3A",x"22",x"15",
    x"C6",x"12",x"D7",x"77",x"86",x"5B",x"BD",x"D6",x"A2",x"DC",x"31",x"BD",x"C4",x"5A",x"86",x"5D",
    x"BD",x"D6",x"A2",x"0F",x"77",x"9D",x"C0",x"8D",x"02",x"20",x"BA",x"BD",x"27",x"C7",x"27",x"B4",
    x"4D",x"10",x"2A",x"E7",x"7A",x"81",x"F8",x"22",x"0B",x"BE",x"27",x"73",x"48",x"1F",x"89",x"3A",
    x"9D",x"C0",x"6E",x"94",x"81",x"FF",x"27",x"04",x"6E",x"9F",x"27",x"7D",x"9D",x"C0",x"81",x"9C",
    x"10",x"27",x"F3",x"77",x"81",x"A1",x"10",x"27",x"FD",x"06",x"81",x"A4",x"10",x"27",x"11",x"13",
    x"81",x"BA",x"25",x"09",x"81",x"C0",x"22",x"05",x"8E",x"CF",x"6A",x"20",x"CF",x"7E",x"27",x"CA",
    x"D6",x"31",x"5C",x"27",x"09",x"C6",x"13",x"7D",x"2C",x"29",x"10",x"26",x"51",x"19",x"5F",x"7E",
    x"B5",x"24",x"42",x"41",x"53",x"44",x"41",x"54",x"42",x"49",x"4E",x"4D",x"41",x"50",x"8E",x"22",
    x"4E",x"6F",x"80",x"CC",x"20",x"13",x"A7",x"80",x"5A",x"26",x"FB",x"39",x"B6",x"27",x"6F",x"BD",
    x"28",x"0C",x"97",x"B2",x"8D",x"E8",x"37",x"24",x"F7",x"22",x"57",x"10",x"BF",x"22",x"58",x"9D",
    x"C6",x"27",x"49",x"BD",x"BF",x"30",x"C1",x"02",x"25",x"18",x"86",x"3A",x"A1",x"01",x"10",x"26",
    x"00",x"83",x"A6",x"81",x"80",x"30",x"25",x"29",x"81",x"09",x"22",x"25",x"8A",x"80",x"97",x"B2",
    x"C0",x"02",x"CE",x"22",x"5A",x"5D",x"27",x"1D",x"A6",x"84",x"81",x"28",x"26",x"17",x"30",x"01",
    x"5A",x"27",x"0E",x"A6",x"80",x"81",x"29",x"27",x"0B",x"A7",x"C0",x"11",x"83",x"22",x"7B",x"25",
    x"EF",x"16",x"00",x"86",x"5A",x"6F",x"C4",x"CE",x"22",x"4F",x"5C",x"5A",x"27",x"46",x"A6",x"80",
    x"81",x"2E",x"27",x"0D",x"11",x"83",x"22",x"57",x"27",x"E7",x"8D",x"21",x"7C",x"22",x"4E",x"20",
    x"EA",x"CE",x"22",x"5A",x"86",x"20",x"A7",x"C2",x"11",x"83",x"22",x"57",x"26",x"F8",x"5A",x"27",
    x"23",x"A6",x"80",x"11",x"83",x"22",x"5A",x"27",x"C8",x"8D",x"02",x"20",x"F1",x"A7",x"C0",x"27",
    x"C0",x"81",x"28",x"27",x"BC",x"81",x"29",x"27",x"B8",x"81",x"3A",x"27",x"B4",x"81",x"2E",x"27",
    x"B0",x"4C",x"27",x"AD",x"39",x"C1",x"05",x"25",x"89",x"A1",x"04",x"26",x"85",x"34",x"14",x"C6",
    x"0F",x"D7",x"B2",x"CE",x"29",x"1A",x"D6",x"B2",x"58",x"EE",x"C5",x"27",x"16",x"AE",x"61",x"C6",
    x"04",x"A6",x"C0",x"A1",x"80",x"26",x"0C",x"5A",x"26",x"F7",x"35",x"14",x"30",x"05",x"C0",x"05",
    x"7E",x"D0",x"F2",x"0A",x"B2",x"2A",x"DC",x"7E",x"D4",x"57",x"C6",x"37",x"0E",x"B7",x"81",x"22",
    x"26",x"21",x"8D",x"06",x"27",x"1D",x"9D",x"BA",x"20",x"19",x"CE",x"D0",x"A2",x"BD",x"D0",x"BC",
    x"C6",x"11",x"D7",x"77",x"7F",x"22",x"4C",x"7F",x"22",x"4D",x"7F",x"28",x"17",x"0E",x"C6",x"9D",
    x"C0",x"26",x"A1",x"7F",x"2C",x"44",x"BD",x"C4",x"CF",x"8D",x"3E",x"73",x"22",x"4D",x"73",x"28",
    x"17",x"0D",x"77",x"27",x"03",x"BD",x"D4",x"1D",x"9E",x"6B",x"7E",x"C4",x"66",x"81",x"4D",x"10",
    x"27",x"01",x"30",x"81",x"50",x"10",x"27",x"00",x"B7",x"8D",x"BF",x"27",x"24",x"9D",x"BA",x"81",
    x"41",x"27",x"CC",x"C6",x"50",x"9D",x"BD",x"26",x"09",x"86",x"FF",x"20",x"17",x"CC",x"0B",x"0D",
    x"DD",x"D9",x"39",x"9E",x"31",x"30",x"01",x"26",x"79",x"0D",x"79",x"27",x"75",x"C6",x"3D",x"0E",
    x"B7",x"8D",x"F6",x"4F",x"97",x"D8",x"BD",x"D2",x"EF",x"96",x"D8",x"4A",x"8D",x"65",x"8D",x"DD",
    x"96",x"21",x"81",x"02",x"22",x"0F",x"5F",x"4A",x"27",x"02",x"86",x"40",x"D3",x"1F",x"80",x"60",
    x"BD",x"D3",x"0B",x"20",x"09",x"DC",x"1F",x"BD",x"D3",x"0B",x"96",x"21",x"8D",x"45",x"4F",x"4C",
    x"34",x"02",x"BD",x"DC",x"19",x"10",x"8E",x"60",x"01",x"20",x"08",x"A6",x"A0",x"8D",x"17",x"30",
    x"1F",x"26",x"F8",x"AE",x"A4",x"26",x"F4",x"35",x"02",x"E6",x"22",x"26",x"E2",x"4F",x"8D",x"06",
    x"4F",x"8D",x"03",x"7E",x"D3",x"4F",x"0D",x"D8",x"27",x"19",x"90",x"D9",x"8D",x"18",x"9B",x"DA",
    x"8D",x"11",x"0A",x"D9",x"26",x"04",x"C6",x"0B",x"D7",x"D9",x"0A",x"DA",x"26",x"04",x"C6",x"0D",
    x"D7",x"DA",x"39",x"7E",x"D6",x"A2",x"CE",x"D8",x"96",x"D6",x"D9",x"A8",x"C5",x"CE",x"D8",x"89",
    x"D6",x"DA",x"A8",x"C5",x"39",x"9D",x"C0",x"CE",x"D0",x"AB",x"BD",x"D1",x"AD",x"7E",x"E4",x"55",
    x"8D",x"F3",x"8D",x"3E",x"CE",x"ED",x"C0",x"BD",x"B0",x"02",x"8D",x"5F",x"8D",x"5B",x"8D",x"0B",
    x"8D",x"15",x"86",x"FF",x"8D",x"57",x"8D",x"51",x"7E",x"D3",x"4A",x"9E",x"45",x"96",x"47",x"97",
    x"DE",x"30",x"02",x"CE",x"D2",x"D3",x"39",x"AD",x"C4",x"A6",x"80",x"BD",x"D6",x"A2",x"31",x"3F",
    x"26",x"F5",x"39",x"8C",x"9F",x"F7",x"23",x"3A",x"34",x"40",x"CE",x"ED",x"1B",x"BD",x"B0",x"02",
    x"35",x"C0",x"BD",x"C1",x"E1",x"86",x"02",x"B7",x"22",x"4C",x"8D",x"03",x"4F",x"20",x"1E",x"BD",
    x"D4",x"1D",x"7D",x"22",x"4D",x"26",x"08",x"B6",x"22",x"19",x"80",x"03",x"B7",x"22",x"B0",x"39",
    x"BD",x"C1",x"64",x"35",x"40",x"34",x"10",x"6E",x"C4",x"4F",x"5F",x"8D",x"00",x"BD",x"D6",x"A2",
    x"1E",x"89",x"39",x"9D",x"C0",x"CE",x"D0",x"A8",x"BD",x"D1",x"AD",x"8D",x"E3",x"8D",x"E1",x"AC",
    x"62",x"10",x"25",x"EC",x"1E",x"8D",x"D9",x"BD",x"C5",x"2B",x"8D",x"B6",x"EC",x"62",x"A3",x"64",
    x"C3",x"00",x"01",x"1F",x"02",x"8D",x"D4",x"EC",x"64",x"8D",x"D0",x"AE",x"64",x"CE",x"D3",x"12",
    x"8D",x"85",x"86",x"FF",x"8D",x"C7",x"8D",x"C1",x"35",x"36",x"8D",x"BF",x"BD",x"DC",x"23",x"D6",
    x"77",x"0F",x"77",x"8E",x"29",x"3A",x"3A",x"BD",x"27",x"EE",x"A6",x"84",x"27",x"16",x"B7",x"22",
    x"B0",x"2B",x"12",x"34",x"10",x"84",x"30",x"B7",x"22",x"4B",x"E6",x"84",x"BD",x"D6",x"BB",x"AD",
    x"98",x"06",x"6F",x"F1",x"39",x"84",x"0F",x"B7",x"22",x"44",x"E6",x"84",x"6F",x"84",x"C5",x"40",
    x"27",x"03",x"BD",x"EA",x"9A",x"CE",x"B6",x"E1",x"7E",x"B0",x"02",x"27",x"0C",x"8D",x"18",x"8D",
    x"BE",x"9D",x"C6",x"27",x"0F",x"8D",x"0E",x"20",x"F6",x"C6",x"11",x"34",x"04",x"8D",x"B2",x"35",
    x"04",x"5A",x"2A",x"F7",x"39",x"9D",x"BA",x"9D",x"C6",x"81",x"23",x"26",x"02",x"9D",x"C0",x"C6",
    x"10",x"BD",x"C1",x"E9",x"D7",x"77",x"26",x"EC",x"C6",x"32",x"0E",x"B7",x"F6",x"22",x"B1",x"4F",
    x"1F",x"01",x"9D",x"C6",x"27",x"03",x"BD",x"C1",x"64",x"BF",x"22",x"47",x"26",x"D6",x"7E",x"BF",
    x"43",x"BD",x"B9",x"06",x"BD",x"BE",x"F5",x"34",x"04",x"8D",x"CA",x"BD",x"D6",x"EB",x"26",x"7A",
    x"9D",x"BA",x"CE",x"D0",x"A5",x"BD",x"D0",x"BC",x"8D",x"D2",x"9D",x"C6",x"26",x"51",x"CC",x"01",
    x"FF",x"FD",x"22",x"4C",x"F7",x"28",x"17",x"35",x"04",x"8D",x"24",x"0F",x"77",x"7C",x"28",x"17",
    x"27",x"3D",x"BD",x"DF",x"39",x"20",x"4D",x"96",x"B2",x"2B",x"06",x"81",x"02",x"10",x"26",x"53",
    x"AD",x"C6",x"11",x"D7",x"77",x"8D",x"03",x"7E",x"D2",x"F2",x"C6",x"49",x"8C",x"C6",x"4F",x"BD",
    x"27",x"EB",x"8D",x"1C",x"B7",x"22",x"4B",x"D6",x"B2",x"2B",x"33",x"BD",x"D6",x"BB",x"27",x"27",
    x"AD",x"98",x"04",x"96",x"B2",x"BA",x"22",x"4B",x"8E",x"29",x"3A",x"D6",x"77",x"A7",x"85",x"39",
    x"86",x"10",x"C1",x"49",x"27",x"F9",x"48",x"C1",x"4F",x"27",x"F4",x"48",x"C1",x"52",x"27",x"EF",
    x"C1",x"44",x"27",x"EB",x"C6",x"33",x"8C",x"C6",x"3C",x"8C",x"C6",x"34",x"0E",x"B7",x"84",x"40",
    x"27",x"13",x"FC",x"22",x"AA",x"F3",x"22",x"47",x"34",x"06",x"25",x"05",x"B3",x"27",x"6D",x"23",
    x"04",x"C6",x"49",x"0E",x"B7",x"BD",x"E7",x"D1",x"CE",x"B4",x"AD",x"BD",x"B0",x"02",x"B6",x"22",
    x"4B",x"85",x"40",x"27",x"05",x"35",x"06",x"FD",x"22",x"AA",x"86",x"80",x"BA",x"22",x"44",x"20",
    x"A4",x"86",x"02",x"B7",x"29",x"50",x"20",x"18",x"CC",x"00",x"FF",x"F7",x"29",x"50",x"20",x"14",
    x"81",x"50",x"10",x"27",x"01",x"AD",x"80",x"4D",x"B7",x"29",x"50",x"26",x"02",x"9D",x"C0",x"4F",
    x"5F",x"FD",x"29",x"51",x"B7",x"29",x"4E",x"F7",x"29",x"4F",x"CE",x"D0",x"A2",x"7D",x"29",x"50",
    x"26",x"03",x"CE",x"D0",x"A8",x"BD",x"D0",x"BC",x"7D",x"29",x"50",x"26",x"0B",x"BD",x"B8",x"E7",
    x"27",x"06",x"BD",x"C1",x"66",x"BF",x"29",x"51",x"BD",x"B8",x"E7",x"27",x"0C",x"C6",x"52",x"9D",
    x"BD",x"BD",x"C5",x"2B",x"86",x"03",x"B7",x"29",x"4E",x"BD",x"D4",x"07",x"7D",x"29",x"50",x"10",
    x"27",x"01",x"12",x"FC",x"22",x"4C",x"27",x"2B",x"5D",x"26",x"06",x"BD",x"D3",x"4F",x"7E",x"D4",
    x"54",x"96",x"B2",x"81",x"02",x"26",x"05",x"7D",x"28",x"17",x"27",x"EF",x"7D",x"29",x"4F",x"26",
    x"03",x"BD",x"B4",x"2E",x"7E",x"B2",x"A8",x"BD",x"D5",x"FA",x"4C",x"97",x"79",x"BD",x"D1",x"FD",
    x"7E",x"D6",x"32",x"7D",x"29",x"4F",x"26",x"D3",x"BD",x"B4",x"2E",x"73",x"29",x"53",x"8D",x"E7",
    x"4D",x"2A",x"07",x"1F",x"01",x"BD",x"D5",x"FA",x"20",x"15",x"6F",x"E2",x"8B",x"60",x"25",x"06",
    x"10",x"83",x"9F",x"FF",x"25",x"04",x"6C",x"E4",x"80",x"40",x"1F",x"01",x"35",x"02",x"4C",x"BD",
    x"B3",x"B9",x"86",x"01",x"BD",x"DC",x"19",x"97",x"6D",x"8E",x"60",x"01",x"9F",x"D6",x"10",x"8E",
    x"00",x"00",x"8D",x"11",x"8D",x"0F",x"D6",x"78",x"26",x"42",x"8D",x"0B",x"26",x"FC",x"10",x"AF",
    x"9F",x"21",x"D6",x"20",x"E7",x"8D",x"00",x"BD",x"D6",x"81",x"D6",x"79",x"27",x"0A",x"90",x"DA",
    x"BD",x"D2",x"86",x"9B",x"D9",x"BD",x"D2",x"72",x"8C",x"9F",x"FC",x"26",x"1A",x"34",x"02",x"DC",
    x"D6",x"FD",x"9F",x"FE",x"CC",x"60",x"01",x"DD",x"D6",x"30",x"AB",x"0C",x"6D",x"96",x"6D",x"BD",
    x"DC",x"19",x"7F",x"60",x"00",x"35",x"02",x"31",x"21",x"A7",x"80",x"39",x"9E",x"D6",x"8D",x"43",
    x"96",x"6D",x"BD",x"B3",x"B9",x"4A",x"27",x"23",x"97",x"70",x"BD",x"DC",x"19",x"10",x"BE",x"9F",
    x"FE",x"CE",x"9F",x"FC",x"8E",x"60",x"03",x"6F",x"A0",x"6F",x"A0",x"34",x"20",x"BD",x"DC",x"32",
    x"0A",x"6D",x"96",x"6D",x"BD",x"DC",x"19",x"A7",x"F1",x"20",x"DA",x"BD",x"D3",x"4F",x"BD",x"B4",
    x"3D",x"77",x"29",x"4E",x"25",x"03",x"BD",x"D3",x"99",x"77",x"29",x"4E",x"10",x"25",x"FA",x"15",
    x"7E",x"B2",x"9B",x"6F",x"80",x"6F",x"80",x"6F",x"84",x"39",x"BD",x"D6",x"81",x"0D",x"78",x"27",
    x"F8",x"C6",x"35",x"0E",x"B7",x"BD",x"C1",x"E1",x"8D",x"2F",x"8D",x"EE",x"34",x"02",x"8D",x"22",
    x"1F",x"02",x"8D",x"1E",x"F3",x"29",x"51",x"FD",x"27",x"A8",x"1F",x"01",x"A6",x"E0",x"26",x"07",
    x"CE",x"D6",x"52",x"8D",x"1F",x"20",x"E3",x"BD",x"D3",x"4F",x"7D",x"29",x"4E",x"27",x"4F",x"7E",
    x"C2",x"0E",x"8D",x"00",x"8D",x"C4",x"1E",x"89",x"39",x"FC",x"22",x"4C",x"83",x"02",x"00",x"27",
    x"F7",x"7E",x"D4",x"FB",x"8D",x"3B",x"D6",x"78",x"26",x"B7",x"AD",x"C4",x"A7",x"80",x"31",x"3F",
    x"26",x"F2",x"39",x"BD",x"D2",x"95",x"BD",x"D4",x"07",x"8D",x"DE",x"CE",x"EB",x"9E",x"BD",x"B0",
    x"02",x"34",x"06",x"8D",x"95",x"8D",x"CB",x"1F",x"02",x"A3",x"E1",x"10",x"24",x"DB",x"8D",x"8D",
    x"C1",x"BD",x"D2",x"BB",x"8D",x"CE",x"CE",x"EB",x"8B",x"8D",x"24",x"BD",x"D3",x"4F",x"7E",x"DC",
    x"23",x"34",x"74",x"BD",x"27",x"F4",x"0F",x"78",x"8D",x"5F",x"2B",x"07",x"8D",x"2D",x"AD",x"98",
    x"08",x"35",x"F4",x"C4",x"0F",x"F7",x"22",x"44",x"CE",x"B6",x"8B",x"8D",x"02",x"35",x"F4",x"7E",
    x"B0",x"02",x"34",x"76",x"BD",x"27",x"F1",x"8D",x"40",x"2B",x"07",x"8D",x"0E",x"AD",x"98",x"0A",
    x"35",x"F6",x"C4",x"0F",x"CE",x"B7",x"D1",x"8D",x"E6",x"35",x"F6",x"C4",x"0F",x"58",x"8E",x"29",
    x"1A",x"AE",x"85",x"39",x"34",x"16",x"BD",x"27",x"F7",x"7F",x"29",x"4D",x"8D",x"1B",x"2B",x"10",
    x"8D",x"E9",x"AD",x"98",x"0C",x"BF",x"2C",x"36",x"FD",x"2C",x"34",x"7D",x"2C",x"37",x"35",x"96",
    x"C4",x"0F",x"CE",x"B8",x"56",x"8D",x"B8",x"20",x"EC",x"D6",x"77",x"8E",x"29",x"3A",x"E6",x"85",
    x"39",x"34",x"14",x"8D",x"F4",x"C4",x"8F",x"35",x"94",x"86",x"20",x"8C",x"86",x"10",x"BD",x"28",
    x"12",x"34",x"16",x"D6",x"77",x"27",x"13",x"8D",x"E2",x"26",x"04",x"C6",x"39",x"0E",x"B7",x"F5",
    x"00",x"40",x"26",x"06",x"E4",x"E4",x"10",x"27",x"FD",x"3A",x"35",x"96",x"8D",x"22",x"BD",x"27",
    x"FA",x"8E",x"29",x"3A",x"6D",x"85",x"10",x"2B",x"13",x"1D",x"96",x"77",x"34",x"02",x"D7",x"77",
    x"8D",x"CA",x"35",x"02",x"97",x"77",x"E6",x"85",x"8D",x"81",x"AD",x"98",x"0E",x"7E",x"BD",x"D4",
    x"BD",x"C1",x"55",x"5A",x"C1",x"0F",x"10",x"22",x"FC",x"6E",x"5C",x"39",x"C6",x"24",x"9D",x"BD",
    x"BD",x"B8",x"DA",x"BD",x"C1",x"4E",x"96",x"77",x"34",x"06",x"0F",x"77",x"9D",x"C6",x"81",x"29",
    x"27",x"03",x"BD",x"D3",x"A5",x"BD",x"B8",x"D7",x"8D",x"92",x"8E",x"23",x"2F",x"E6",x"61",x"27",
    x"0B",x"BD",x"D6",x"81",x"BD",x"CD",x"78",x"A7",x"80",x"5A",x"26",x"F5",x"35",x"06",x"97",x"77",
    x"7E",x"BF",x"68",x"9D",x"C6",x"81",x"28",x"26",x"0C",x"BD",x"B8",x"D3",x"BD",x"C1",x"55",x"5D",
    x"27",x"03",x"8D",x"AF",x"21",x"5F",x"96",x"77",x"34",x"02",x"D7",x"77",x"BD",x"D6",x"F9",x"BD",
    x"D6",x"C4",x"35",x"02",x"97",x"77",x"F6",x"2C",x"36",x"7E",x"BD",x"D6",x"BD",x"D1",x"AA",x"BD",
    x"B8",x"E7",x"BD",x"C5",x"A0",x"8D",x"43",x"BD",x"D4",x"07",x"FC",x"22",x"4C",x"10",x"26",x"FC",
    x"93",x"BD",x"D5",x"17",x"4D",x"2A",x"03",x"BD",x"D5",x"FA",x"8E",x"29",x"56",x"10",x"8E",x"00",
    x"00",x"BD",x"D5",x"75",x"BD",x"D5",x"75",x"0D",x"78",x"26",x"11",x"BD",x"D5",x"77",x"26",x"FB",
    x"FC",x"29",x"58",x"DD",x"33",x"1F",x"20",x"BD",x"B2",x"FA",x"20",x"DE",x"BD",x"D3",x"4F",x"B6",
    x"2C",x"3C",x"4C",x"10",x"27",x"DC",x"29",x"7E",x"B6",x"AB",x"8E",x"2A",x"5E",x"CE",x"00",x"00",
    x"A6",x"84",x"44",x"44",x"25",x"02",x"EF",x"01",x"44",x"25",x"02",x"EF",x"03",x"30",x"07",x"8C",
    x"2B",x"14",x"26",x"EC",x"9E",x"1B",x"33",x"84",x"20",x"1E",x"10",x"AE",x"84",x"A6",x"02",x"BD",
    x"DC",x"14",x"F1",x"2B",x"D2",x"25",x"0F",x"22",x"06",x"10",x"BC",x"2B",x"D0",x"25",x"07",x"E6",
    x"03",x"10",x"AF",x"C1",x"ED",x"C1",x"30",x"04",x"9C",x"1D",x"26",x"DE",x"DF",x"1D",x"BE",x"2B",
    x"D0",x"B6",x"2B",x"D2",x"9F",x"25",x"97",x"27",x"39",x"8D",x"AF",x"9D",x"C6",x"26",x"10",x"9E",
    x"25",x"96",x"27",x"BF",x"2B",x"D0",x"B7",x"2B",x"D2",x"39",x"BD",x"B8",x"E7",x"27",x"F0",x"9E",
    x"C7",x"A6",x"80",x"27",x"11",x"81",x"3A",x"27",x"0D",x"81",x"2C",x"27",x"09",x"81",x"28",x"26",
    x"F0",x"BD",x"BC",x"25",x"20",x"E4",x"BD",x"BB",x"96",x"4D",x"26",x"09",x"4C",x"90",x"05",x"D6",
    x"05",x"EA",x"86",x"E7",x"86",x"BD",x"DC",x"23",x"20",x"D0",x"86",x"1E",x"D7",x"BA",x"87",x"99",
    x"26",x"64",x"87",x"23",x"34",x"58",x"86",x"80",x"19",x"56",x"AA",x"80",x"76",x"22",x"F1",x"82",
    x"38",x"AA",x"BD",x"C1",x"55",x"C1",x"10",x"10",x"24",x"E6",x"98",x"8E",x"1F",x"FF",x"10",x"8E",
    x"00",x"00",x"1F",x"98",x"8D",x"52",x"1F",x"10",x"88",x"10",x"85",x"10",x"27",x"03",x"53",x"88",
    x"EF",x"DD",x"50",x"39",x"C6",x"0F",x"BD",x"C1",x"E9",x"34",x"04",x"8E",x"1F",x"FF",x"4F",x"5F",
    x"34",x"06",x"BD",x"B8",x"E7",x"27",x"14",x"BD",x"C1",x"66",x"DC",x"50",x"2A",x"02",x"43",x"53",
    x"ED",x"E4",x"81",x"10",x"10",x"24",x"E6",x"5B",x"8E",x"10",x"00",x"34",x"10",x"BD",x"B8",x"E7",
    x"27",x"12",x"A6",x"E4",x"84",x"EF",x"A7",x"E4",x"BD",x"E0",x"F5",x"5D",x"26",x"06",x"C6",x"10",
    x"EA",x"62",x"E7",x"62",x"35",x"30",x"35",x"02",x"3F",x"BC",x"BD",x"27",x"FD",x"7D",x"23",x"01",
    x"26",x"0B",x"C6",x"05",x"F7",x"23",x"01",x"3F",x"0C",x"27",x"02",x"8D",x"36",x"7D",x"2B",x"34",
    x"27",x"A1",x"7D",x"2C",x"29",x"26",x"9C",x"BD",x"C9",x"A7",x"8E",x"2B",x"37",x"20",x"47",x"BD",
    x"27",x"FD",x"3F",x"0C",x"27",x"8D",x"34",x"04",x"3F",x"0A",x"5D",x"27",x"14",x"C1",x"03",x"10",
    x"27",x"DB",x"D3",x"C1",x"02",x"26",x"07",x"3F",x"0A",x"5D",x"27",x"FB",x"20",x"EF",x"F7",x"2B",
    x"69",x"35",x"84",x"34",x"14",x"8D",x"DF",x"27",x"1B",x"7D",x"2C",x"29",x"26",x"16",x"8E",x"2B",
    x"3D",x"F6",x"2B",x"69",x"30",x"04",x"E1",x"84",x"26",x"FA",x"8C",x"2B",x"69",x"27",x"05",x"7F",
    x"2B",x"69",x"20",x"02",x"35",x"94",x"10",x"DE",x"75",x"96",x"31",x"4C",x"27",x"19",x"D6",x"1A",
    x"DE",x"C7",x"A6",x"03",x"34",x"01",x"84",x"7F",x"97",x"1A",x"BD",x"DC",x"19",x"AE",x"01",x"9F",
    x"C7",x"35",x"01",x"2A",x"02",x"8D",x"03",x"7E",x"D0",x"05",x"10",x"9E",x"31",x"86",x"BC",x"34",
    x"66",x"20",x"F4",x"C6",x"18",x"8C",x"C6",x"07",x"8C",x"C6",x"0C",x"3F",x"82",x"F6",x"20",x"1B",
    x"20",x"16",x"8D",x"02",x"20",x"12",x"BD",x"C1",x"55",x"C1",x"01",x"10",x"22",x"E5",x"84",x"1F",
    x"98",x"3F",x"9C",x"8D",x"F1",x"25",x"17",x"5F",x"7E",x"BD",x"D4",x"BD",x"C1",x"55",x"C1",x"01",
    x"10",x"22",x"E5",x"6F",x"5C",x"34",x"04",x"BD",x"DA",x"DD",x"E4",x"E0",x"27",x"E9",x"C6",x"FF",
    x"20",x"E6",x"3F",x"16",x"20",x"DF",x"26",x"0E",x"8E",x"2B",x"D7",x"CC",x"FF",x"40",x"A7",x"80",
    x"5A",x"26",x"FB",x"39",x"9D",x"BA",x"C6",x"07",x"BD",x"C1",x"E9",x"34",x"04",x"C6",x"3B",x"9D",
    x"BD",x"27",x"3C",x"81",x"2C",x"27",x"38",x"BD",x"E2",x"2B",x"27",x"3C",x"81",x"2C",x"27",x"38",
    x"34",x"30",x"C6",x"C8",x"9D",x"BD",x"BD",x"E2",x"2B",x"E6",x"64",x"86",x"08",x"3D",x"CE",x"2B",
    x"D7",x"33",x"CB",x"8D",x"0D",x"32",x"62",x"1F",x"21",x"8D",x"07",x"32",x"63",x"9D",x"C6",x"26",
    x"C3",x"39",x"EC",x"62",x"AC",x"62",x"24",x"02",x"1E",x"01",x"ED",x"C1",x"AF",x"42",x"39",x"8E",
    x"FF",x"FF",x"1F",x"12",x"34",x"30",x"20",x"D1",x"BD",x"E2",x"53",x"1F",x"10",x"5A",x"86",x"08",
    x"3D",x"1F",x"01",x"1F",x"20",x"86",x"08",x"3D",x"1F",x"02",x"34",x"30",x"30",x"07",x"31",x"27",
    x"20",x"B7",x"81",x"B8",x"10",x"26",x"DC",x"EE",x"9D",x"C0",x"8D",x"65",x"25",x"1D",x"CE",x"2B",
    x"D7",x"5F",x"5C",x"AC",x"C4",x"25",x"0E",x"10",x"AC",x"42",x"25",x"09",x"AC",x"44",x"22",x"05",
    x"10",x"AC",x"46",x"23",x"07",x"33",x"48",x"C1",x"08",x"26",x"E7",x"5F",x"D7",x"51",x"7E",x"B7",
    x"6B",x"9D",x"C0",x"BD",x"D9",x"2F",x"8D",x"45",x"27",x"F9",x"8D",x"49",x"20",x"06",x"9D",x"C0",
    x"8D",x"27",x"8D",x"2F",x"34",x"30",x"8D",x"1B",x"35",x"40",x"8D",x"06",x"9D",x"BA",x"8D",x"13",
    x"35",x"40",x"DF",x"50",x"C6",x"02",x"D7",x"05",x"BD",x"B0",x"27",x"9E",x"45",x"BD",x"B0",x"33",
    x"7E",x"DC",x"23",x"BD",x"BB",x"96",x"96",x"05",x"39",x"BD",x"D9",x"2F",x"3F",x"16",x"24",x"F9",
    x"39",x"8D",x"F6",x"3F",x"18",x"24",x"05",x"8E",x"FF",x"FF",x"1F",x"12",x"39",x"5F",x"3F",x"3E",
    x"26",x"01",x"5C",x"59",x"39",x"3F",x"40",x"20",x"EC",x"9D",x"C0",x"C6",x"99",x"9D",x"BD",x"BD",
    x"B8",x"DA",x"F6",x"2C",x"17",x"10",x"27",x"E4",x"4A",x"5A",x"BD",x"C1",x"E9",x"86",x"08",x"97",
    x"F4",x"3D",x"F3",x"20",x"70",x"DD",x"F2",x"BD",x"B8",x"D7",x"C6",x"D4",x"9D",x"BD",x"8C",x"9D",
    x"BA",x"BD",x"C1",x"4E",x"34",x"04",x"0A",x"F4",x"26",x"F5",x"86",x"08",x"9E",x"F2",x"35",x"04",
    x"E7",x"80",x"4A",x"26",x"F9",x"39",x"22",x"41",x"55",x"54",x"4F",x"2E",x"42",x"41",x"54",x"00",
    x"10",x"DE",x"28",x"CE",x"B1",x"36",x"BD",x"B0",x"02",x"F6",x"29",x"53",x"27",x"03",x"BD",x"B4",
    x"2E",x"BD",x"B4",x"3F",x"BD",x"D3",x"99",x"8D",x"06",x"BD",x"28",x"0F",x"7E",x"B2",x"9B",x"BD",
    x"E3",x"BE",x"BD",x"C3",x"53",x"1B",x"66",x"1B",x"44",x"1B",x"56",x"0C",x"11",x"00",x"86",x"04",
    x"B7",x"2C",x"4A",x"8E",x"23",x"00",x"BF",x"20",x"61",x"B7",x"20",x"63",x"39",x"CC",x"C6",x"21",
    x"1F",x"9B",x"7F",x"2D",x"1A",x"B1",x"23",x"00",x"27",x"B6",x"10",x"CE",x"5F",x"FF",x"CE",x"B1",
    x"41",x"BD",x"B0",x"02",x"03",x"31",x"10",x"FF",x"2C",x"4B",x"BD",x"DD",x"37",x"86",x"02",x"7D",
    x"20",x"80",x"27",x"10",x"CE",x"BD",x"D0",x"BD",x"B0",x"02",x"86",x"02",x"8E",x"01",x"00",x"BD",
    x"E9",x"8D",x"86",x"80",x"B7",x"27",x"6F",x"8D",x"A6",x"BD",x"B4",x"2E",x"BD",x"C3",x"53",x"42",
    x"41",x"53",x"49",x"43",x"20",x"31",x"32",x"38",x"20",x"56",x"31",x"2E",x"30",x"20",x"28",x"63",
    x"29",x"20",x"4D",x"69",x"63",x"72",x"6F",x"73",x"6F",x"66",x"74",x"20",x"31",x"39",x"38",x"36",
    x"0D",x"0A",x"00",x"8E",x"DB",x"26",x"9F",x"C7",x"7D",x"20",x"80",x"27",x"06",x"7E",x"D4",x"91",
    x"BD",x"B4",x"2E",x"CE",x"D3",x"BA",x"BD",x"B0",x"02",x"BD",x"BF",x"89",x"BD",x"C3",x"34",x"BD",
    x"C3",x"53",x"20",x"62",x"79",x"74",x"65",x"73",x"20",x"66",x"72",x"65",x"65",x"00",x"7E",x"B2",
    x"9B",x"A6",x"80",x"A7",x"C0",x"5A",x"26",x"F9",x"39",x"4F",x"34",x"40",x"A7",x"80",x"AC",x"E4",
    x"23",x"FA",x"35",x"C0",x"1F",x"89",x"D0",x"8A",x"39",x"A7",x"E2",x"27",x"04",x"9B",x"8A",x"8D",
    x"06",x"35",x"82",x"96",x"1A",x"9B",x"8A",x"B7",x"A7",x"E5",x"97",x"8B",x"39",x"10",x"9E",x"6E",
    x"9E",x"6B",x"1F",x"40",x"83",x"00",x"14",x"34",x"47",x"1A",x"50",x"96",x"70",x"91",x"6D",x"26",
    x"06",x"8D",x"D6",x"8D",x"3A",x"20",x"1C",x"DE",x"1D",x"96",x"70",x"8D",x"CC",x"20",x"04",x"A6",
    x"A0",x"A7",x"C0",x"10",x"AC",x"63",x"24",x"09",x"11",x"A3",x"61",x"26",x"F2",x"8D",x"0B",x"20",
    x"E6",x"8D",x"07",x"9F",x"6B",x"10",x"9F",x"6E",x"35",x"C7",x"34",x"40",x"96",x"6D",x"8D",x"A9",
    x"DE",x"1D",x"20",x"04",x"A6",x"C0",x"A7",x"80",x"11",x"A3",x"E4",x"26",x"F7",x"35",x"C0",x"34",
    x"20",x"AC",x"E1",x"25",x"17",x"1F",x"30",x"34",x"20",x"A3",x"E4",x"30",x"8B",x"34",x"50",x"20",
    x"04",x"A6",x"C2",x"A7",x"82",x"11",x"A3",x"64",x"26",x"F7",x"35",x"F0",x"34",x"40",x"20",x"04",
    x"A6",x"A0",x"A7",x"80",x"10",x"AC",x"E4",x"25",x"F7",x"35",x"C0",x"4B",x"59",x"42",x"44",x"DC",
    x"BB",x"DC",x"C9",x"DC",x"C2",x"DC",x"DC",x"DD",x"0D",x"DC",x"CA",x"81",x"10",x"27",x"0A",x"7E",
    x"D4",x"54",x"3F",x"0A",x"5D",x"27",x"FB",x"1F",x"98",x"39",x"5F",x"39",x"53",x"43",x"52",x"4E",
    x"DD",x"08",x"DD",x"0C",x"DC",x"C2",x"DC",x"DC",x"DD",x"0D",x"D4",x"54",x"81",x"0D",x"26",x"08",
    x"7D",x"20",x"2C",x"2A",x"03",x"BD",x"D9",x"A3",x"F6",x"20",x"2A",x"C4",x"01",x"27",x"15",x"34",
    x"02",x"B6",x"20",x"1B",x"4A",x"2B",x"05",x"8E",x"22",x"00",x"6F",x"86",x"35",x"02",x"81",x"0A",
    x"26",x"02",x"8D",x"00",x"1F",x"89",x"3F",x"82",x"81",x"20",x"26",x"B3",x"39",x"B6",x"20",x"1C",
    x"4A",x"BD",x"E2",x"6E",x"1F",x"01",x"86",x"0D",x"C0",x"28",x"27",x"02",x"C6",x"27",x"CB",x"1A",
    x"39",x"03",x"06",x"07",x"08",x"0A",x"0C",x"0E",x"0F",x"C0",x"00",x"40",x"80",x"B7",x"20",x"82",
    x"3F",x"C2",x"B7",x"20",x"42",x"3F",x"A4",x"8E",x"DD",x"2D",x"BF",x"2C",x"1D",x"30",x"05",x"BF",
    x"2C",x"24",x"39",x"9D",x"C0",x"8E",x"2C",x"1F",x"A6",x"84",x"34",x"02",x"26",x"02",x"8D",x"2C",
    x"17",x"00",x"88",x"86",x"02",x"8D",x"34",x"A6",x"E0",x"27",x"27",x"39",x"4C",x"50",x"52",x"54",
    x"DD",x"6C",x"DD",x"82",x"D4",x"54",x"DD",x"95",x"DD",x"D1",x"D4",x"54",x"8D",x"9A",x"8E",x"2C",
    x"1F",x"6D",x"84",x"10",x"26",x"01",x"D8",x"CE",x"22",x"5A",x"8D",x"6D",x"63",x"84",x"86",x"04",
    x"20",x"09",x"8E",x"2C",x"1F",x"8D",x"54",x"6F",x"84",x"86",x"10",x"AD",x"98",x"05",x"24",x"90",
    x"8D",x"F5",x"7E",x"DF",x"4C",x"8E",x"2C",x"1F",x"6D",x"04",x"26",x"04",x"81",x"16",x"26",x"06",
    x"63",x"04",x"39",x"8E",x"2C",x"18",x"81",x"0D",x"26",x"04",x"6F",x"01",x"20",x"18",x"81",x"20",
    x"25",x"14",x"E6",x"02",x"27",x"10",x"E1",x"01",x"22",x"08",x"34",x"02",x"8D",x"21",x"35",x"02",
    x"6F",x"01",x"6C",x"01",x"27",x"F4",x"1F",x"89",x"86",x"01",x"20",x"BF",x"8E",x"2C",x"18",x"20",
    x"03",x"8E",x"2C",x"1F",x"86",x"0D",x"E6",x"03",x"AE",x"01",x"39",x"6D",x"01",x"27",x"39",x"6F",
    x"01",x"86",x"0D",x"8D",x"E1",x"86",x"0A",x"20",x"DD",x"6F",x"01",x"C6",x"28",x"A6",x"C4",x"27",
    x"18",x"10",x"9E",x"C7",x"34",x"30",x"DF",x"C7",x"9D",x"C6",x"BD",x"B7",x"8E",x"DC",x"33",x"4D",
    x"10",x"26",x"E1",x"3F",x"35",x"30",x"10",x"9F",x"C7",x"E7",x"02",x"4F",x"8B",x"0D",x"25",x"04",
    x"A1",x"02",x"23",x"F8",x"80",x"1A",x"A7",x"03",x"39",x"43",x"4F",x"4D",x"4D",x"DE",x"29",x"DE",
    x"79",x"DE",x"8C",x"DD",x"A3",x"DD",x"CC",x"DC",x"CA",x"8E",x"2C",x"18",x"CE",x"22",x"5A",x"A5",
    x"84",x"10",x"26",x"01",x"1A",x"AA",x"84",x"E6",x"84",x"A7",x"84",x"5D",x"26",x"DA",x"C6",x"04",
    x"A6",x"C4",x"27",x"06",x"33",x"41",x"80",x"31",x"1F",x"89",x"C1",x"08",x"22",x"28",x"10",x"8E",
    x"DD",x"21",x"E6",x"A5",x"F7",x"20",x"85",x"C6",x"40",x"A6",x"C4",x"27",x"0E",x"33",x"41",x"80",
    x"35",x"2D",x"13",x"81",x"03",x"22",x"0F",x"31",x"28",x"E6",x"A6",x"EA",x"04",x"F7",x"20",x"84",
    x"17",x"FF",x"76",x"16",x"FF",x"08",x"7E",x"BF",x"43",x"8E",x"2C",x"18",x"43",x"A4",x"84",x"A7",
    x"84",x"10",x"27",x"FF",x"00",x"84",x"20",x"10",x"27",x"FF",x"50",x"39",x"4F",x"C6",x"02",x"F7",
    x"20",x"82",x"3F",x"42",x"25",x"02",x"1F",x"98",x"39",x"43",x"41",x"53",x"53",x"DE",x"D4",x"DF",
    x"27",x"DE",x"CC",x"DF",x"5B",x"DE",x"A9",x"DE",x"C3",x"73",x"29",x"4D",x"CC",x"01",x"00",x"8E",
    x"00",x"00",x"39",x"D6",x"B4",x"E0",x"3F",x"A6",x"AB",x"6A",x"3F",x"26",x"16",x"34",x"02",x"8D",
    x"7E",x"35",x"82",x"BD",x"DF",x"53",x"26",x"01",x"43",x"1E",x"89",x"39",x"BD",x"DF",x"53",x"26",
    x"E2",x"03",x"78",x"39",x"0D",x"B5",x"26",x"77",x"81",x"10",x"10",x"27",x"00",x"93",x"8E",x"22",
    x"4E",x"6D",x"80",x"10",x"27",x"F2",x"B3",x"CE",x"28",x"1B",x"C6",x"0B",x"BD",x"DC",x"01",x"B6",
    x"20",x"79",x"E6",x"84",x"C0",x"31",x"26",x"02",x"8A",x"04",x"5A",x"26",x"02",x"84",x"FC",x"B7",
    x"20",x"79",x"FC",x"22",x"4C",x"ED",x"C1",x"B6",x"28",x"17",x"A7",x"C0",x"C6",x"0E",x"E7",x"51",
    x"86",x"02",x"97",x"B5",x"0F",x"B3",x"F7",x"28",x"18",x"BD",x"DF",x"C2",x"B6",x"28",x"17",x"B7",
    x"28",x"18",x"8D",x"2F",x"6F",x"3F",x"39",x"0D",x"B5",x"27",x"13",x"81",x"20",x"26",x"0A",x"8D",
    x"22",x"27",x"02",x"8D",x"53",x"C6",x"FF",x"8D",x"51",x"BD",x"DF",x"E1",x"0F",x"B5",x"39",x"8D",
    x"69",x"27",x"07",x"2B",x"04",x"8D",x"0C",x"27",x"F6",x"39",x"8D",x"ED",x"C6",x"35",x"8C",x"C6",
    x"3B",x"0E",x"B7",x"10",x"8E",x"28",x"1B",x"4F",x"E6",x"3F",x"39",x"34",x"02",x"8D",x"F4",x"CB",
    x"02",x"26",x"04",x"8D",x"23",x"C6",x"02",x"5A",x"E7",x"3F",x"31",x"AB",x"35",x"02",x"A7",x"3F",
    x"39",x"BD",x"DF",x"F7",x"8D",x"AC",x"EC",x"2B",x"FD",x"22",x"4C",x"A6",x"2D",x"B7",x"28",x"17",
    x"B7",x"28",x"18",x"8D",x"BA",x"0C",x"B5",x"39",x"C6",x"01",x"D7",x"B3",x"8D",x"34",x"20",x"92",
    x"86",x"02",x"CE",x"D0",x"A2",x"BD",x"D0",x"BF",x"96",x"B2",x"81",x"02",x"10",x"26",x"DF",x"A3",
    x"8D",x"CF",x"0D",x"B3",x"2B",x"93",x"8D",x"97",x"20",x"F8",x"8D",x"41",x"10",x"8E",x"28",x"1A",
    x"3F",x"20",x"4D",x"26",x"95",x"A6",x"A0",x"80",x"02",x"97",x"B4",x"A7",x"3F",x"8D",x"1D",x"D7",
    x"B3",x"39",x"8D",x"29",x"8D",x"8D",x"30",x"A4",x"5D",x"27",x"05",x"AB",x"80",x"5A",x"26",x"FB",
    x"40",x"A7",x"84",x"6C",x"A2",x"6C",x"A4",x"4F",x"D6",x"B3",x"3F",x"20",x"7D",x"28",x"18",x"27",
    x"15",x"4F",x"B7",x"2D",x"1A",x"3F",x"22",x"24",x"0D",x"C6",x"3C",x"0E",x"B7",x"96",x"B5",x"8A",
    x"01",x"7D",x"2D",x"1A",x"27",x"EC",x"39",x"96",x"31",x"4C",x"B7",x"28",x"19",x"8E",x"E0",x"59",
    x"8D",x"23",x"7F",x"28",x"18",x"8D",x"A3",x"26",x"F9",x"8D",x"D6",x"8E",x"22",x"4E",x"6D",x"80",
    x"27",x"0B",x"C6",x"0B",x"A6",x"80",x"A1",x"A0",x"26",x"13",x"5A",x"26",x"F7",x"8E",x"E0",x"67",
    x"8D",x"21",x"8E",x"E0",x"64",x"7D",x"28",x"19",x"26",x"CC",x"7E",x"C3",x"4E",x"8E",x"E0",x"6F",
    x"8D",x"11",x"20",x"C9",x"1F",x"89",x"9D",x"C0",x"C1",x"96",x"27",x"B1",x"C1",x"C3",x"27",x"A1",
    x"7E",x"B8",x"F4",x"8D",x"E0",x"7D",x"28",x"19",x"26",x"DE",x"8E",x"28",x"1B",x"C6",x"08",x"8D",
    x"05",x"BD",x"C3",x"47",x"C6",x"03",x"7E",x"C3",x"39",x"0D",x"0A",x"53",x"65",x"61",x"72",x"63",
    x"68",x"69",x"6E",x"67",x"0D",x"0A",x"00",x"46",x"6F",x"75",x"6E",x"64",x"3A",x"20",x"00",x"53",
    x"6B",x"69",x"70",x"3A",x"20",x"00",x"8E",x"2D",x"1B",x"9F",x"E0",x"8E",x"29",x"5B",x"31",x"89",
    x"00",x"FF",x"BD",x"D6",x"F1",x"26",x"0A",x"0F",x"78",x"CE",x"DB",x"23",x"BD",x"B0",x"02",x"20",
    x"23",x"BD",x"D6",x"81",x"0D",x"78",x"26",x"13",x"81",x"0D",x"27",x"0F",x"81",x"16",x"27",x"04",
    x"81",x"20",x"25",x"ED",x"A7",x"80",x"8C",x"2A",x"5A",x"25",x"E6",x"BD",x"D6",x"F1",x"10",x"2B",
    x"0A",x"FC",x"6F",x"84",x"8E",x"29",x"5A",x"39",x"F6",x"20",x"1C",x"81",x"2C",x"27",x"07",x"BD",
    x"E2",x"6E",x"5A",x"8D",x"32",x"5C",x"B6",x"20",x"1B",x"34",x"06",x"BD",x"B8",x"E7",x"27",x"06",
    x"C6",x"18",x"8D",x"23",x"E7",x"E4",x"9D",x"C6",x"27",x"0B",x"8D",x"17",x"27",x"03",x"C6",x"14",
    x"8C",x"C6",x"11",x"8D",x"0C",x"C6",x"1F",x"8D",x"08",x"35",x"04",x"8D",x"02",x"35",x"04",x"CB",
    x"40",x"3F",x"82",x"9D",x"BA",x"C6",x"01",x"7E",x"C1",x"E9",x"C6",x"02",x"8D",x"02",x"C6",x"01",
    x"9D",x"C6",x"27",x"1F",x"81",x"2C",x"27",x"19",x"34",x"04",x"53",x"F4",x"20",x"2A",x"34",x"04",
    x"8D",x"E3",x"27",x"02",x"6F",x"61",x"35",x"04",x"EA",x"E0",x"F7",x"20",x"2A",x"9D",x"C6",x"27",
    x"02",x"0E",x"BA",x"39",x"C6",x"02",x"20",x"CF",x"F6",x"20",x"1E",x"81",x"2C",x"27",x"04",x"C6",
    x"18",x"8D",x"C4",x"34",x"04",x"F6",x"20",x"20",x"BD",x"B8",x"E7",x"27",x"04",x"C6",x"18",x"8D",
    x"B6",x"E1",x"E4",x"10",x"25",x"DD",x"FC",x"CE",x"DD",x"24",x"BD",x"B0",x"02",x"35",x"04",x"CE",
    x"DD",x"21",x"BD",x"B0",x"02",x"BD",x"B8",x"E7",x"27",x"18",x"C6",x"07",x"BD",x"C1",x"E9",x"4F",
    x"54",x"D7",x"A0",x"C6",x"74",x"24",x"02",x"43",x"5C",x"B7",x"22",x"88",x"17",x"00",x"8B",x"BD",
    x"E2",x"CD",x"BD",x"B8",x"E7",x"27",x"07",x"8D",x"AB",x"CB",x"78",x"17",x"00",x"7C",x"BD",x"B8",
    x"E7",x"27",x"A0",x"C6",x"0B",x"BD",x"C1",x"E9",x"CB",x"7C",x"17",x"00",x"6D",x"BD",x"E2",x"CD",
    x"7E",x"E3",x"BE",x"9D",x"C0",x"81",x"AB",x"10",x"27",x"FB",x"A8",x"C6",x"5F",x"F7",x"2B",x"14",
    x"9D",x"C6",x"27",x"11",x"81",x"2C",x"27",x"0D",x"17",x"00",x"6A",x"F7",x"2C",x"4A",x"BD",x"E2",
    x"C7",x"CA",x"40",x"8D",x"48",x"BD",x"B8",x"E7",x"27",x"06",x"8D",x"59",x"CA",x"50",x"8D",x"3D",
    x"7D",x"2B",x"14",x"27",x"0E",x"BD",x"B8",x"E7",x"27",x"09",x"8D",x"49",x"CA",x"60",x"8D",x"2A",
    x"73",x"2B",x"14",x"BD",x"B8",x"E7",x"27",x"14",x"BD",x"E0",x"F5",x"C6",x"7B",x"8D",x"1E",x"F6",
    x"20",x"2B",x"54",x"54",x"54",x"54",x"F7",x"2C",x"4A",x"BD",x"E2",x"C7",x"7D",x"2B",x"14",x"27",
    x"23",x"9D",x"C6",x"27",x"1F",x"BD",x"E0",x"F3",x"CB",x"76",x"7F",x"2B",x"14",x"34",x"04",x"C6",
    x"1B",x"8D",x"0F",x"7D",x"2B",x"14",x"27",x"08",x"C6",x"23",x"8D",x"06",x"C6",x"20",x"8D",x"02",
    x"35",x"04",x"3F",x"82",x"39",x"C6",x"0F",x"7E",x"C1",x"E9",x"8D",x"0F",x"3F",x"14",x"7E",x"BD",
    x"D4",x"8D",x"08",x"8D",x"2E",x"CE",x"D3",x"35",x"7E",x"B0",x"02",x"9D",x"C6",x"81",x"C6",x"34",
    x"01",x"26",x"02",x"9D",x"C0",x"BD",x"B8",x"DA",x"BD",x"BA",x"A2",x"34",x"10",x"BD",x"BA",x"A0",
    x"31",x"84",x"35",x"10",x"35",x"01",x"26",x"08",x"DC",x"A1",x"30",x"8B",x"DC",x"A3",x"31",x"AB",
    x"7E",x"B8",x"D7",x"8D",x"19",x"4F",x"34",x"06",x"30",x"01",x"27",x"06",x"AC",x"E4",x"22",x"02",
    x"AF",x"E4",x"10",x"8C",x"00",x"18",x"23",x"04",x"10",x"8E",x"00",x"18",x"35",x"90",x"F6",x"20",
    x"77",x"2B",x"0A",x"C4",x"40",x"26",x"03",x"C6",x"28",x"39",x"C6",x"14",x"39",x"C6",x"50",x"39",
    x"BD",x"E3",x"25",x"8D",x"1A",x"CE",x"E1",x"4F",x"20",x"0B",x"81",x"FF",x"10",x"27",x"EA",x"4C",
    x"8D",x"6E",x"CE",x"E4",x"41",x"7D",x"20",x"36",x"10",x"26",x"00",x"D2",x"7E",x"B0",x"02",x"7F",
    x"20",x"36",x"F6",x"20",x"2A",x"D7",x"66",x"F6",x"2C",x"4A",x"9D",x"C6",x"27",x"19",x"81",x"3B",
    x"27",x"15",x"81",x"2C",x"26",x"26",x"BD",x"BA",x"A0",x"DC",x"50",x"10",x"83",x"FF",x"F0",x"2D",
    x"7F",x"10",x"83",x"00",x"0F",x"2E",x"79",x"D1",x"9F",x"27",x"B4",x"D7",x"9F",x"CE",x"E3",x"16",
    x"7E",x"B0",x"02",x"34",x"76",x"F6",x"2C",x"4A",x"8D",x"ED",x"35",x"F6",x"BD",x"E3",x"EB",x"C1",
    x"20",x"25",x"5D",x"F7",x"20",x"36",x"B6",x"20",x"2A",x"84",x"FC",x"B7",x"20",x"2A",x"9E",x"A1",
    x"10",x"9E",x"A3",x"8D",x"23",x"8D",x"31",x"9D",x"C6",x"27",x"32",x"9D",x"BA",x"7E",x"E1",x"9C",
    x"81",x"C8",x"27",x"02",x"8D",x"1F",x"C6",x"C8",x"9D",x"BD",x"BD",x"E2",x"2B",x"34",x"30",x"8D",
    x"8E",x"35",x"30",x"7D",x"20",x"36",x"27",x"15",x"7E",x"E2",x"53",x"0F",x"EF",x"81",x"46",x"26",
    x"0C",x"03",x"EF",x"0E",x"C0",x"BD",x"E2",x"2B",x"9F",x"A1",x"10",x"9F",x"A3",x"39",x"8D",x"EB",
    x"8D",x"F3",x"81",x"2C",x"27",x"0D",x"BD",x"C1",x"4E",x"D7",x"F1",x"BD",x"C1",x"60",x"20",x"08",
    x"7E",x"BF",x"43",x"BD",x"C1",x"60",x"D7",x"F1",x"D7",x"F0",x"BD",x"E4",x"06",x"0F",x"F2",x"9D",
    x"C6",x"81",x"3B",x"26",x"16",x"9D",x"C0",x"03",x"F2",x"BD",x"BA",x"AD",x"8E",x"21",x"F3",x"BD",
    x"B0",x"33",x"BD",x"BA",x"AB",x"8E",x"21",x"F7",x"BD",x"B0",x"33",x"CE",x"DF",x"96",x"BD",x"B0",
    x"02",x"96",x"66",x"B7",x"20",x"2A",x"39",x"8D",x"A2",x"8D",x"85",x"CE",x"E7",x"56",x"20",x"EE",
    x"BD",x"E2",x"2B",x"10",x"AF",x"E3",x"2D",x"B8",x"AF",x"E3",x"2D",x"B4",x"C6",x"C8",x"9D",x"BD",
    x"BD",x"E2",x"2B",x"10",x"8C",x"00",x"C8",x"24",x"A7",x"8D",x"1C",x"34",x"06",x"AC",x"E1",x"24",
    x"9F",x"AC",x"E4",x"25",x"9B",x"10",x"AC",x"62",x"25",x"96",x"9F",x"A9",x"10",x"9F",x"AB",x"35",
    x"30",x"9F",x"A5",x"10",x"9F",x"A7",x"39",x"BD",x"E2",x"6E",x"86",x"08",x"3D",x"39",x"8D",x"F7",
    x"5A",x"DD",x"A9",x"4F",x"5F",x"DD",x"A5",x"DD",x"A7",x"CC",x"00",x"C7",x"DD",x"AB",x"39",x"8D",
    x"1A",x"C1",x"20",x"25",x"D3",x"BE",x"20",x"73",x"5D",x"2A",x"05",x"BE",x"20",x"70",x"C0",x"60",
    x"C0",x"1F",x"86",x"08",x"3D",x"30",x"8B",x"BF",x"22",x"7D",x"39",x"BD",x"B9",x"06",x"BD",x"B9",
    x"45",x"10",x"26",x"DD",x"60",x"7E",x"BE",x"F5",x"BD",x"E3",x"25",x"8D",x"09",x"BD",x"EC",x"3D",
    x"CE",x"E7",x"B2",x"16",x"FF",x"68",x"BD",x"E2",x"9F",x"7D",x"20",x"36",x"27",x"DC",x"7E",x"B8",
    x"F4",x"8D",x"32",x"34",x"06",x"9D",x"C6",x"81",x"2C",x"26",x"08",x"8D",x"1E",x"1F",x"98",x"C6",
    x"18",x"20",x"06",x"C6",x"C8",x"9D",x"BD",x"8D",x"1C",x"34",x"06",x"BD",x"E2",x"D3",x"8D",x"25",
    x"35",x"30",x"CE",x"EB",x"66",x"BD",x"B0",x"02",x"7E",x"DC",x"23",x"BD",x"E2",x"6E",x"C1",x"14",
    x"26",x"02",x"C6",x"50",x"39",x"BD",x"E2",x"2B",x"8D",x"F1",x"BD",x"E2",x"55",x"34",x"30",x"A6",
    x"61",x"E6",x"63",x"35",x"B0",x"9D",x"BA",x"C6",x"80",x"D7",x"04",x"BD",x"BB",x"12",x"27",x"AE",
    x"D6",x"05",x"C1",x"82",x"10",x"26",x"DA",x"D5",x"BD",x"BD",x"5A",x"E1",x"80",x"26",x"9F",x"5A",
    x"26",x"9C",x"EC",x"E4",x"DD",x"6B",x"EC",x"02",x"DD",x"6E",x"A6",x"04",x"97",x"70",x"BD",x"BC",
    x"C1",x"9F",x"45",x"97",x"47",x"8D",x"B1",x"BD",x"C5",x"2B",x"96",x"47",x"7E",x"DC",x"19",x"BD",
    x"BF",x"30",x"31",x"84",x"96",x"51",x"CE",x"DE",x"A7",x"BD",x"B0",x"02",x"BD",x"B8",x"E7",x"26",
    x"EE",x"39",x"30",x"64",x"97",x"E7",x"A6",x"84",x"C6",x"0C",x"81",x"EF",x"27",x"06",x"81",x"81",
    x"26",x"1F",x"C6",x"19",x"91",x"E7",x"26",x"0F",x"A6",x"03",x"DE",x"48",x"27",x"0C",x"11",x"A3",
    x"01",x"26",x"04",x"91",x"4A",x"27",x"09",x"3A",x"20",x"DC",x"EE",x"01",x"DF",x"48",x"97",x"4A",
    x"4F",x"39",x"BD",x"B6",x"EC",x"9F",x"E2",x"96",x"1A",x"97",x"E4",x"9E",x"31",x"9F",x"DF",x"96",
    x"8B",x"97",x"E1",x"39",x"35",x"20",x"CE",x"21",x"E5",x"C6",x"06",x"A6",x"C2",x"34",x"02",x"5A",
    x"26",x"F9",x"6E",x"A4",x"35",x"20",x"9E",x"31",x"96",x"1A",x"34",x"12",x"9E",x"C7",x"34",x"10",
    x"6E",x"A4",x"BD",x"B7",x"B3",x"27",x"05",x"BD",x"B9",x"42",x"24",x"03",x"7E",x"BF",x"3D",x"8E",
    x"21",x"67",x"BD",x"B0",x"33",x"BD",x"DC",x"23",x"32",x"62",x"8D",x"B6",x"30",x"E4",x"86",x"81",
    x"8D",x"82",x"26",x"11",x"3A",x"EC",x"1D",x"93",x"E2",x"26",x"F3",x"A6",x"1F",x"90",x"E4",x"26",
    x"ED",x"32",x"84",x"9F",x"75",x"C6",x"0D",x"BD",x"B1",x"E1",x"8D",x"A8",x"C6",x"BB",x"BD",x"B7",
    x"BE",x"D6",x"56",x"CA",x"7F",x"D4",x"4F",x"9E",x"50",x"96",x"4E",x"34",x"16",x"8E",x"00",x"01",
    x"9F",x"50",x"BD",x"B9",x"42",x"22",x"09",x"8E",x"D0",x"EE",x"CE",x"C1",x"84",x"BD",x"B0",x"02",
    x"9D",x"C6",x"81",x"C6",x"26",x"08",x"9D",x"C0",x"BD",x"B7",x"C0",x"BD",x"DC",x"23",x"CE",x"C2",
    x"56",x"BD",x"B0",x"02",x"34",x"04",x"DE",x"50",x"9E",x"4E",x"96",x"05",x"34",x"52",x"BD",x"C5",
    x"2B",x"CC",x"81",x"82",x"BD",x"E6",x"7A",x"BD",x"E4",x"F4",x"D6",x"4A",x"34",x"04",x"9E",x"48",
    x"C6",x"81",x"34",x"17",x"86",x"4F",x"97",x"71",x"8E",x"00",x"00",x"9F",x"48",x"9E",x"C7",x"9F",
    x"E5",x"9D",x"C6",x"27",x"07",x"BD",x"BB",x"96",x"9F",x"48",x"97",x"4A",x"86",x"81",x"BD",x"E4",
    x"A2",x"27",x"04",x"C6",x"01",x"0E",x"B7",x"96",x"4A",x"BD",x"DC",x"27",x"32",x"84",x"A6",x"66",
    x"91",x"1A",x"26",x"EF",x"AE",x"64",x"9C",x"E5",x"26",x"E9",x"A6",x"69",x"97",x"05",x"81",x"02",
    x"27",x"31",x"CE",x"D3",x"94",x"BD",x"B0",x"02",x"E0",x"6E",x"27",x"0F",x"EE",x"E8",x"13",x"A6",
    x"E8",x"15",x"E6",x"E8",x"18",x"AE",x"E8",x"16",x"7E",x"E6",x"6E",x"32",x"E8",x"19",x"30",x"E4",
    x"9F",x"75",x"BD",x"DC",x"23",x"9D",x"C6",x"81",x"2C",x"10",x"26",x"EA",x"08",x"9D",x"C0",x"0F",
    x"71",x"8D",x"98",x"9E",x"48",x"96",x"71",x"26",x"0A",x"EC",x"84",x"E3",x"6C",x"28",x"06",x"C6",
    x"06",x"0E",x"B7",x"DC",x"67",x"ED",x"84",x"A3",x"E8",x"11",x"27",x"BC",x"2C",x"04",x"C6",x"FF",
    x"20",x"B6",x"C6",x"01",x"20",x"B2",x"32",x"62",x"BD",x"E4",x"D2",x"CC",x"EF",x"F0",x"8D",x"4A",
    x"96",x"1A",x"97",x"4A",x"9E",x"C7",x"9F",x"48",x"30",x"E4",x"86",x"EF",x"BD",x"E4",x"A4",x"26",
    x"05",x"32",x"85",x"10",x"DF",x"75",x"C6",x"06",x"BD",x"B1",x"E1",x"BD",x"E4",x"E4",x"BD",x"E4",
    x"F4",x"C6",x"EF",x"34",x"07",x"9E",x"C7",x"9F",x"48",x"96",x"1A",x"97",x"4A",x"86",x"EF",x"BD",
    x"E4",x"A2",x"26",x"45",x"32",x"84",x"EE",x"66",x"AE",x"69",x"E6",x"6B",x"A6",x"68",x"DF",x"31",
    x"9F",x"C7",x"D7",x"1A",x"BD",x"DC",x"27",x"7E",x"D0",x"05",x"34",x"06",x"5F",x"5C",x"9D",x"C6",
    x"20",x"02",x"9D",x"C0",x"27",x"08",x"81",x"8F",x"27",x"25",x"81",x"C4",x"26",x"F4",x"4D",x"26",
    x"1E",x"9E",x"C7",x"30",x"01",x"BD",x"CF",x"EC",x"26",x"13",x"9E",x"DF",x"9F",x"31",x"C6",x"17",
    x"35",x"02",x"81",x"81",x"27",x"05",x"C6",x"19",x"8C",x"C6",x"1A",x"0E",x"B7",x"DF",x"31",x"9D",
    x"C0",x"A1",x"E4",x"27",x"C8",x"A1",x"61",x"26",x"C5",x"5A",x"26",x"04",x"9D",x"C0",x"35",x"86",
    x"9D",x"C0",x"27",x"CA",x"34",x"04",x"BD",x"BB",x"7C",x"35",x"04",x"BD",x"DC",x"23",x"9D",x"C6",
    x"27",x"BC",x"81",x"2C",x"27",x"E3",x"7E",x"B8",x"F4",x"C6",x"01",x"9D",x"C6",x"27",x"03",x"BD",
    x"C1",x"4E",x"D7",x"D6",x"26",x"01",x"39",x"C6",x"02",x"32",x"E5",x"A6",x"E4",x"33",x"64",x"31",
    x"E8",x"16",x"C6",x"19",x"81",x"81",x"27",x"0E",x"33",x"61",x"31",x"69",x"C6",x"0C",x"81",x"EF",
    x"27",x"04",x"C6",x"18",x"0E",x"B7",x"96",x"1A",x"9E",x"C7",x"A1",x"42",x"22",x"DB",x"26",x"04",
    x"AC",x"C4",x"22",x"D5",x"A1",x"22",x"25",x"D1",x"26",x"04",x"AC",x"A4",x"25",x"CB",x"0A",x"D6",
    x"26",x"C7",x"A6",x"42",x"97",x"1A",x"BD",x"DC",x"23",x"AE",x"C4",x"9F",x"C7",x"AE",x"43",x"9F",
    x"31",x"32",x"E5",x"C1",x"EF",x"27",x"02",x"9D",x"C6",x"10",x"27",x"E8",x"C8",x"BD",x"BB",x"7C",
    x"7E",x"E5",x"EE",x"CE",x"22",x"4F",x"C6",x"13",x"20",x"05",x"CE",x"20",x"48",x"C6",x"09",x"35",
    x"20",x"33",x"C5",x"A6",x"C2",x"34",x"02",x"5A",x"26",x"F9",x"6E",x"A4",x"CE",x"20",x"48",x"C6",
    x"09",x"35",x"20",x"35",x"02",x"A7",x"C0",x"5A",x"26",x"F9",x"6E",x"A4",x"8D",x"28",x"8D",x"DA",
    x"BD",x"BF",x"2E",x"8D",x"E7",x"BD",x"BE",x"75",x"F1",x"22",x"B1",x"25",x"03",x"F6",x"22",x"B1",
    x"4F",x"30",x"CB",x"F0",x"22",x"B1",x"50",x"27",x"05",x"A7",x"80",x"5A",x"26",x"FB",x"C6",x"08",
    x"CE",x"B2",x"E7",x"7E",x"B0",x"02",x"8D",x"42",x"34",x"04",x"BD",x"C1",x"60",x"34",x"04",x"BD",
    x"C1",x"60",x"5A",x"C1",x"10",x"10",x"24",x"D7",x"9A",x"5C",x"F7",x"20",x"4C",x"35",x"06",x"B7",
    x"20",x"4B",x"F7",x"20",x"49",x"39",x"BD",x"B8",x"DA",x"8D",x"DB",x"BD",x"B8",x"D7",x"CE",x"23",
    x"2F",x"C6",x"02",x"8D",x"CB",x"F6",x"22",x"B1",x"7E",x"BF",x"68",x"CE",x"E8",x"5A",x"BD",x"D0",
    x"BC",x"D6",x"B2",x"C8",x"80",x"2A",x"06",x"7E",x"D4",x"57",x"BD",x"C1",x"4E",x"7D",x"20",x"80",
    x"27",x"F5",x"F7",x"20",x"49",x"C1",x"04",x"22",x"EE",x"39",x"80",x"C3",x"27",x"08",x"81",x"D3",
    x"10",x"26",x"D1",x"00",x"86",x"80",x"97",x"8D",x"0E",x"C0",x"86",x"FF",x"97",x"B2",x"BD",x"D0",
    x"BF",x"D6",x"B2",x"2A",x"04",x"8D",x"CA",x"CA",x"80",x"F7",x"27",x"6F",x"39",x"BD",x"C1",x"55",
    x"8D",x"CB",x"0C",x"89",x"CE",x"B3",x"6A",x"7E",x"B0",x"02",x"0D",x"77",x"26",x"EE",x"C6",x"7B",
    x"7E",x"E1",x"FA",x"80",x"50",x"34",x"01",x"26",x"02",x"9D",x"C0",x"8D",x"9E",x"35",x"01",x"26",
    x"0A",x"CC",x"11",x"03",x"97",x"77",x"D7",x"B2",x"BD",x"D4",x"1D",x"8D",x"DD",x"F6",x"22",x"B1",
    x"8E",x"E9",x"49",x"5C",x"26",x"02",x"30",x"04",x"C6",x"04",x"BD",x"C3",x"39",x"BD",x"C3",x"53",
    x"6C",x"65",x"20",x"64",x"65",x"6E",x"73",x"69",x"74",x"79",x"20",x"20",x"20",x"00",x"B6",x"20",
    x"49",x"8B",x"30",x"BD",x"D6",x"A2",x"86",x"3A",x"BD",x"D6",x"A2",x"0C",x"89",x"8D",x"AB",x"CE",
    x"B4",x"16",x"8D",x"A3",x"8D",x"A4",x"BD",x"C3",x"34",x"BD",x"C3",x"53",x"20",x"44",x"53",x"4B",
    x"46",x"20",x"3D",x"20",x"00",x"8D",x"93",x"8D",x"8B",x"8D",x"8F",x"BD",x"E9",x"36",x"BD",x"C4",
    x"5F",x"8D",x"87",x"BD",x"C2",x"DD",x"BD",x"C4",x"5F",x"BD",x"C2",x"DD",x"8E",x"22",x"4F",x"A6",
    x"80",x"81",x"20",x"26",x"02",x"6F",x"1F",x"8C",x"22",x"5A",x"26",x"F3",x"CE",x"B3",x"AB",x"20",
    x"03",x"CE",x"B3",x"A0",x"BD",x"B0",x"02",x"96",x"8E",x"10",x"27",x"EA",x"92",x"BD",x"D9",x"2F",
    x"9E",x"8F",x"C6",x"08",x"8D",x"4A",x"C6",x"09",x"8D",x"49",x"C6",x"03",x"8D",x"42",x"C6",x"0D",
    x"8D",x"41",x"86",x"2A",x"E6",x"84",x"C1",x"09",x"22",x"05",x"CE",x"E9",x"3F",x"A6",x"C5",x"8D",
    x"3E",x"A6",x"01",x"8B",x"42",x"8D",x"38",x"8D",x"4D",x"30",x"05",x"6D",x"84",x"2F",x"09",x"C6",
    x"15",x"8D",x"20",x"C6",x"08",x"8D",x"19",x"8C",x"30",x"08",x"6D",x"84",x"2F",x"0A",x"C6",x"1E",
    x"8D",x"11",x"8D",x"22",x"8D",x"20",x"8D",x"24",x"BD",x"C4",x"5F",x"BD",x"C2",x"DD",x"20",x"A1",
    x"7E",x"C3",x"39",x"BD",x"D6",x"C4",x"F0",x"2C",x"36",x"8D",x"06",x"5A",x"26",x"FB",x"39",x"8D",
    x"02",x"86",x"20",x"7E",x"D6",x"A2",x"8D",x"04",x"86",x"2D",x"20",x"F7",x"E6",x"80",x"C1",x"09",
    x"22",x"02",x"8D",x"ED",x"4F",x"8C",x"DC",x"50",x"34",x"10",x"BD",x"C4",x"5A",x"35",x"90",x"42",
    x"44",x"4D",x"41",x"34",x"35",x"36",x"37",x"38",x"39",x"53",x"69",x"6E",x"67",x"44",x"6F",x"75",
    x"62",x"FC",x"27",x"6D",x"93",x"87",x"34",x"06",x"D6",x"95",x"34",x"04",x"9D",x"C6",x"81",x"2C",
    x"8D",x"21",x"BD",x"B8",x"E7",x"27",x"05",x"BD",x"C1",x"66",x"AF",x"61",x"BD",x"D3",x"99",x"35",
    x"12",x"8D",x"1A",x"F6",x"2C",x"4D",x"BD",x"B8",x"E7",x"27",x"05",x"C6",x"19",x"BD",x"C1",x"E9",
    x"7E",x"B5",x"5A",x"27",x"07",x"C6",x"0F",x"BD",x"C1",x"E9",x"E7",x"62",x"39",x"4C",x"1F",x"89",
    x"34",x"16",x"EC",x"62",x"D3",x"87",x"10",x"25",x"C8",x"62",x"ED",x"62",x"C3",x"01",x"1B",x"25",
    x"F5",x"6A",x"E4",x"26",x"F7",x"C3",x"00",x"04",x"C4",x"FC",x"1F",x"03",x"BD",x"B1",x"E5",x"DF",
    x"1B",x"9E",x"87",x"BF",x"22",x"AA",x"BD",x"DC",x"09",x"35",x"16",x"CE",x"B2",x"BF",x"7E",x"B0",
    x"02",x"BD",x"E7",x"CB",x"BD",x"C5",x"2B",x"CE",x"B4",x"7F",x"20",x"20",x"BD",x"E7",x"DA",x"86",
    x"07",x"34",x"06",x"BD",x"B8",x"E7",x"8D",x"AB",x"BD",x"D3",x"99",x"BD",x"B8",x"E7",x"BD",x"D0",
    x"BC",x"35",x"06",x"B7",x"20",x"4D",x"F7",x"20",x"49",x"CE",x"B8",x"61",x"20",x"5E",x"BD",x"E7",
    x"CB",x"34",x"04",x"BD",x"E7",x"43",x"8D",x"1B",x"BD",x"E7",x"CB",x"E1",x"E8",x"13",x"10",x"26",
    x"D5",x"41",x"BD",x"E7",x"43",x"30",x"E8",x"13",x"31",x"E4",x"CE",x"B8",x"8D",x"8D",x"3D",x"32",
    x"E8",x"27",x"39",x"C6",x"41",x"9D",x"BD",x"C6",x"53",x"0E",x"BD",x"BD",x"D7",x"40",x"8D",x"1E",
    x"CE",x"B8",x"B9",x"20",x"27",x"BD",x"D3",x"A7",x"0F",x"77",x"8D",x"07",x"C5",x"40",x"26",x"14",
    x"7E",x"D4",x"54",x"8E",x"29",x"3A",x"E6",x"85",x"26",x"D8",x"C6",x"39",x"0E",x"B7",x"8D",x"F3",
    x"10",x"2A",x"D4",x"FF",x"C4",x"0F",x"39",x"8D",x"F5",x"CE",x"B8",x"C4",x"7E",x"B0",x"02",x"35",
    x"20",x"CE",x"B4",x"64",x"8D",x"F6",x"EE",x"0B",x"EC",x"09",x"30",x"CB",x"34",x"10",x"34",x"46",
    x"6E",x"A4",x"8D",x"C1",x"8D",x"E9",x"35",x"06",x"9D",x"C6",x"26",x"02",x"35",x"D0",x"BD",x"C1",
    x"60",x"35",x"10",x"4F",x"33",x"8B",x"11",x"A3",x"E4",x"23",x"04",x"C6",x"43",x"0E",x"B7",x"34",
    x"54",x"8D",x"90",x"BD",x"BB",x"96",x"BD",x"BF",x"38",x"35",x"04",x"E7",x"84",x"35",x"06",x"D3",
    x"17",x"93",x"87",x"ED",x"01",x"BD",x"DC",x"23",x"20",x"CE",x"F6",x"22",x"44",x"8D",x"B0",x"DE",
    x"1B",x"20",x"39",x"E6",x"43",x"C5",x"01",x"27",x"31",x"A6",x"42",x"BD",x"DC",x"27",x"AE",x"C4",
    x"E6",x"80",x"3A",x"6D",x"43",x"2A",x"21",x"E6",x"80",x"58",x"3A",x"10",x"AE",x"03",x"A6",x"02",
    x"AE",x"84",x"30",x"1D",x"8C",x"60",x"00",x"24",x"08",x"30",x"89",x"3F",x"F8",x"4A",x"BD",x"DC",
    x"19",x"8D",x"44",x"31",x"3F",x"26",x"EB",x"8C",x"8D",x"3D",x"33",x"44",x"11",x"93",x"1D",x"26",
    x"C2",x"BD",x"DC",x"23",x"D6",x"95",x"34",x"04",x"CE",x"B4",x"64",x"BD",x"B0",x"02",x"A6",x"84",
    x"81",x"40",x"26",x"0B",x"EC",x"0B",x"10",x"A3",x"65",x"25",x"04",x"A3",x"61",x"ED",x"0B",x"35",
    x"04",x"5A",x"2A",x"E2",x"35",x"70",x"20",x"04",x"A6",x"C0",x"A7",x"A0",x"11",x"B3",x"22",x"AA",
    x"26",x"F6",x"10",x"BF",x"22",x"AA",x"39",x"34",x"02",x"EC",x"01",x"93",x"17",x"25",x"12",x"D3",
    x"87",x"10",x"A3",x"65",x"25",x"0B",x"10",x"A3",x"67",x"25",x"08",x"EC",x"01",x"A3",x"63",x"ED",
    x"01",x"35",x"82",x"6F",x"84",x"6F",x"01",x"6F",x"02",x"35",x"82",x"8E",x"29",x"5B",x"C6",x"2C",
    x"D7",x"00",x"BD",x"B9",x"45",x"27",x"02",x"C6",x"20",x"8D",x"73",x"81",x"20",x"27",x"FA",x"81",
    x"22",x"26",x"0A",x"C1",x"2C",x"26",x"06",x"1F",x"89",x"D7",x"00",x"20",x"22",x"C1",x"22",x"27",
    x"11",x"81",x"0D",x"26",x"0D",x"8C",x"29",x"5B",x"27",x"44",x"A6",x"1F",x"81",x"0A",x"26",x"3E",
    x"86",x"0D",x"4D",x"27",x"17",x"91",x"00",x"27",x"1D",x"34",x"04",x"A1",x"E0",x"27",x"17",x"A7",
    x"80",x"8C",x"2A",x"5A",x"26",x"06",x"8D",x"41",x"26",x"06",x"20",x"1E",x"8D",x"3B",x"27",x"CD",
    x"6F",x"84",x"8E",x"29",x"5A",x"39",x"81",x"22",x"27",x"04",x"81",x"20",x"26",x"F2",x"8D",x"29",
    x"26",x"EE",x"81",x"20",x"27",x"F8",x"81",x"2C",x"27",x"E6",x"81",x"0D",x"26",x"08",x"8D",x"19",
    x"26",x"DE",x"81",x"0A",x"27",x"DA",x"CE",x"B8",x"DC",x"BD",x"B0",x"02",x"20",x"D2",x"8D",x"09",
    x"27",x"0C",x"C6",x"36",x"8C",x"C6",x"45",x"0E",x"B7",x"BD",x"D6",x"81",x"0D",x"78",x"39",x"39",
    x"C6",x"5F",x"F7",x"22",x"49",x"81",x"28",x"10",x"27",x"F8",x"36",x"BD",x"EA",x"25",x"F7",x"22",
    x"44",x"8E",x"00",x"00",x"9D",x"C6",x"27",x"07",x"BD",x"C1",x"64",x"9E",x"50",x"27",x"D6",x"CE",
    x"B8",x"FA",x"20",x"09",x"BD",x"D7",x"40",x"BD",x"EA",x"3E",x"CE",x"BA",x"EE",x"7E",x"B0",x"02",
    x"BD",x"E7",x"CB",x"34",x"04",x"BD",x"E7",x"43",x"BD",x"D3",x"99",x"9D",x"C6",x"27",x"17",x"C6",
    x"BB",x"9D",x"BD",x"BD",x"E7",x"CB",x"34",x"04",x"BD",x"E7",x"43",x"30",x"E8",x"14",x"31",x"E4",
    x"8D",x"13",x"32",x"E8",x"28",x"39",x"30",x"E4",x"31",x"E4",x"8D",x"09",x"CE",x"BC",x"7E",x"8D",
    x"1E",x"32",x"E8",x"14",x"39",x"CE",x"BB",x"8E",x"8D",x"C3",x"7E",x"DC",x"23",x"34",x"10",x"9E",
    x"1D",x"9F",x"6B",x"30",x"E8",x"80",x"9F",x"6E",x"35",x"90",x"8E",x"EC",x"FC",x"8D",x"0A",x"8E",
    x"EC",x"F0",x"8D",x"05",x"0D",x"9D",x"26",x"F2",x"39",x"34",x"50",x"BD",x"C3",x"53",x"0C",x"50",
    x"6C",x"65",x"61",x"73",x"65",x"20",x"69",x"6E",x"73",x"65",x"72",x"74",x"20",x"00",x"35",x"10",
    x"BD",x"C3",x"4E",x"BD",x"C3",x"53",x"20",x"64",x"69",x"73",x"6B",x"0D",x"0A",x"26",x"20",x"70",
    x"72",x"65",x"73",x"73",x"20",x"27",x"45",x"4E",x"54",x"52",x"45",x"45",x"27",x"07",x"00",x"3F",
    x"0A",x"C1",x"0D",x"26",x"FA",x"EE",x"E4",x"8D",x"9F",x"35",x"C0",x"BD",x"E7",x"DA",x"34",x"04",
    x"9D",x"C6",x"27",x"07",x"C6",x"BB",x"9D",x"BD",x"BD",x"E7",x"DA",x"35",x"02",x"CE",x"BC",x"AA",
    x"8D",x"86",x"CE",x"BC",x"84",x"0D",x"9D",x"26",x"96",x"39",x"F6",x"27",x"6F",x"9D",x"C6",x"27",
    x"05",x"BD",x"C1",x"4E",x"C8",x"80",x"D7",x"B2",x"BD",x"E7",x"D1",x"C6",x"11",x"34",x"04",x"8E",
    x"29",x"3A",x"E6",x"85",x"2A",x"14",x"C4",x"0F",x"CE",x"B4",x"64",x"BD",x"B0",x"02",x"E6",x"01",
    x"F1",x"20",x"49",x"26",x"05",x"E6",x"E4",x"BD",x"D3",x"51",x"35",x"04",x"5A",x"26",x"DE",x"39",
    x"64",x"65",x"73",x"74",x"69",x"6E",x"61",x"74",x"69",x"6F",x"6E",x"00",x"73",x"6F",x"75",x"72",
    x"63",x"65",x"00",x"8D",x"26",x"26",x"05",x"C6",x"04",x"BD",x"BB",x"BD",x"34",x"12",x"9E",x"C7",
    x"34",x"10",x"BD",x"DC",x"23",x"BD",x"B6",x"E4",x"1F",x"10",x"A3",x"E4",x"35",x"10",x"CE",x"23",
    x"2F",x"D7",x"51",x"BD",x"DC",x"01",x"35",x"42",x"7E",x"B7",x"DC",x"C6",x"BD",x"9D",x"BD",x"86",
    x"40",x"97",x"04",x"7E",x"BB",x"12",x"8D",x"F3",x"26",x"04",x"C6",x"12",x"0E",x"B7",x"4F",x"D6",
    x"05",x"34",x"06",x"BD",x"B8",x"29",x"BD",x"BF",x"4A",x"6F",x"E2",x"30",x"62",x"E6",x"84",x"C1",
    x"28",x"10",x"26",x"00",x"83",x"30",x"01",x"9F",x"73",x"BD",x"B8",x"DA",x"8D",x"52",x"BD",x"BB",
    x"96",x"34",x"12",x"D6",x"05",x"34",x"04",x"BD",x"DC",x"23",x"8D",x"44",x"34",x"06",x"BD",x"B9",
    x"06",x"35",x"10",x"9F",x"73",x"A6",x"E4",x"BD",x"B0",x"27",x"35",x"26",x"81",x"03",x"26",x"17",
    x"4F",x"34",x"12",x"33",x"E4",x"9E",x"2A",x"34",x"10",x"10",x"DF",x"2A",x"34",x"24",x"BD",x"B7",
    x"DC",x"86",x"03",x"34",x"02",x"20",x"0B",x"40",x"32",x"E6",x"40",x"30",x"E4",x"34",x"26",x"BD",
    x"B0",x"33",x"9D",x"C6",x"81",x"29",x"27",x"11",x"9D",x"BA",x"8D",x"04",x"9D",x"BA",x"20",x"AE",
    x"9E",x"73",x"DC",x"C7",x"DD",x"73",x"9F",x"C7",x"39",x"9D",x"C0",x"8D",x"F3",x"BD",x"B8",x"D7",
    x"30",x"E4",x"E6",x"80",x"27",x"16",x"A6",x"80",x"BD",x"DC",x"27",x"EE",x"81",x"C1",x"03",x"26",
    x"02",x"30",x"02",x"BD",x"BD",x"C4",x"20",x"EA",x"9F",x"73",x"8D",x"D4",x"C6",x"D4",x"9D",x"BD",
    x"9E",x"73",x"34",x"10",x"BD",x"B9",x"06",x"35",x"10",x"9F",x"C7",x"30",x"E4",x"E6",x"80",x"27",
    x"16",x"A6",x"80",x"BD",x"DC",x"27",x"EE",x"81",x"C1",x"03",x"26",x"06",x"10",x"AE",x"81",x"10",
    x"9F",x"2A",x"BD",x"DC",x"01",x"20",x"E6",x"E6",x"80",x"4F",x"32",x"8B",x"BD",x"DC",x"23",x"32",
    x"61",x"35",x"02",x"84",x"0F",x"7E",x"B0",x"27",x"8D",x"63",x"E6",x"2E",x"20",x"0A",x"8D",x"5D",
    x"E6",x"2C",x"20",x"04",x"8D",x"57",x"E6",x"2D",x"7E",x"BD",x"D6",x"8D",x"50",x"E6",x"2F",x"C5",
    x"01",x"27",x"09",x"7E",x"D9",x"DE",x"8D",x"45",x"A6",x"2F",x"2B",x"F7",x"7E",x"D9",x"C7",x"BD",
    x"BA",x"A2",x"CE",x"EA",x"2A",x"8D",x"36",x"BD",x"E2",x"D3",x"10",x"8E",x"23",x"2F",x"BD",x"B0",
    x"02",x"8D",x"1A",x"4F",x"33",x"84",x"7E",x"B7",x"DC",x"8D",x"05",x"CE",x"E9",x"4C",x"20",x"E5",
    x"80",x"BB",x"34",x"02",x"26",x"02",x"9D",x"C0",x"BD",x"BA",x"A2",x"35",x"82",x"F6",x"2B",x"15",
    x"10",x"2B",x"D0",x"CF",x"58",x"FB",x"2B",x"15",x"8E",x"2B",x"16",x"3A",x"39",x"34",x"56",x"8D",
    x"EC",x"BD",x"B8",x"29",x"10",x"8E",x"23",x"2F",x"35",x"D6",x"8D",x"D4",x"CE",x"E9",x"45",x"20",
    x"B4",x"8D",x"CD",x"CE",x"E9",x"37",x"20",x"AD",x"8D",x"05",x"CE",x"E9",x"18",x"20",x"A6",x"BD",
    x"BA",x"A2",x"4F",x"30",x"84",x"27",x"01",x"43",x"39",x"81",x"2C",x"27",x"07",x"8D",x"F0",x"CE",
    x"E9",x"2B",x"8D",x"91",x"BD",x"B8",x"E7",x"27",x"EF",x"8D",x"E4",x"CE",x"E9",x"1E",x"20",x"85",
    x"C6",x"09",x"BD",x"C1",x"E9",x"F7",x"2B",x"15",x"8D",x"69",x"9D",x"C6",x"27",x"DA",x"8D",x"AD",
    x"AE",x"26",x"10",x"AE",x"29",x"34",x"30",x"9D",x"BA",x"81",x"2C",x"27",x"05",x"BD",x"BA",x"A2",
    x"AF",x"E4",x"BD",x"B8",x"E7",x"27",x"05",x"BD",x"BA",x"A2",x"AF",x"62",x"8D",x"8F",x"35",x"50",
    x"AF",x"26",x"EF",x"29",x"CE",x"EA",x"62",x"8D",x"37",x"9D",x"C6",x"27",x"AB",x"10",x"8E",x"23",
    x"2F",x"A6",x"2F",x"34",x"22",x"4F",x"CE",x"E9",x"2B",x"BD",x"B0",x"02",x"C6",x"FF",x"D7",x"51",
    x"BD",x"BF",x"4A",x"BD",x"BF",x"2E",x"31",x"84",x"30",x"E8",x"11",x"CE",x"EA",x"D5",x"BD",x"B0",
    x"02",x"4F",x"CB",x"10",x"10",x"25",x"D0",x"18",x"BD",x"BE",x"CC",x"35",x"22",x"CE",x"E9",x"2B",
    x"16",x"FF",x"14",x"BD",x"EE",x"6D",x"6D",x"84",x"26",x"09",x"C6",x"1B",x"D7",x"51",x"CE",x"EA",
    x"B0",x"20",x"ED",x"39",x"9D",x"C0",x"17",x"FF",x"34",x"AE",x"A4",x"10",x"AE",x"22",x"7E",x"DA",
    x"A4",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7E",x"D0",x"BC",x"7E",x"BE",x"1E",x"7E",x"B7",x"D8",
    x"7E",x"BB",x"12",x"7E",x"BC",x"C1",x"7E",x"DC",x"23",x"7E",x"BA",x"A0",x"7E",x"C1",x"64",x"7E",
    x"BA",x"AB",x"7E",x"BF",x"2E",x"7E",x"B9",x"06",x"7E",x"BB",x"96",x"7E",x"B0",x"1D",x"DB",x"6D");

  CONSTANT ROM_MO6_0 : arr8 := (
    x"A6",x"E4",x"84",x"F0",x"A7",x"E4",x"1F",x"8A",x"86",x"20",x"1F",x"8B",x"E6",x"F8",x"0A",x"C4",
    x"7F",x"CE",x"A7",x"C0",x"9E",x"6A",x"EC",x"85",x"85",x"F0",x"26",x"0F",x"8E",x"F0",x"37",x"8A",
    x"F0",x"34",x"16",x"A6",x"C4",x"8A",x"20",x"A7",x"C4",x"20",x"07",x"8E",x"F0",x"43",x"8A",x"00",
    x"34",x"16",x"EC",x"65",x"AE",x"68",x"39",x"34",x"01",x"B6",x"A7",x"C0",x"8A",x"20",x"B7",x"A7",
    x"C0",x"35",x"01",x"1F",x"A8",x"84",x"8F",x"AA",x"E4",x"A7",x"E4",x"AE",x"6A",x"E6",x"80",x"2B",
    x"03",x"AF",x"6A",x"3B",x"35",x"7F",x"32",x"62",x"39",x"01",x"9F",x"F6",x"C7",x"FC",x"09",x"FC",
    x"00",x"FB",x"99",x"F5",x"08",x"02",x"C3",x"06",x"69",x"04",x"A3",x"04",x"C1",x"04",x"E7",x"07",
    x"FA",x"08",x"24",x"FE",x"60",x"0A",x"C1",x"09",x"5A",x"03",x"44",x"04",x"64",x"09",x"D2",x"A0",
    x"04",x"A0",x"07",x"A0",x"0A",x"A0",x"1C",x"A0",x"19",x"A0",x"16",x"A0",x"22",x"A0",x"0D",x"A0",
    x"1F",x"A0",x"10",x"A0",x"13",x"0C",x"71",x"0C",x"E2",x"0C",x"F7",x"0A",x"E7",x"6E",x"9F",x"20",
    x"5E",x"6E",x"9F",x"20",x"67",x"3B",x"3B",x"3B",x"3B",x"3B",x"3B",x"3B",x"3B",x"3B",x"C1",x"05",
    x"23",x"05",x"C1",x"FB",x"24",x"01",x"58",x"1D",x"39",x"C6",x"20",x"1F",x"9B",x"CE",x"A7",x"C0",
    x"96",x"79",x"48",x"2A",x"06",x"A6",x"4E",x"85",x"C0",x"26",x"79",x"A6",x"43",x"85",x"01",x"27",
    x"03",x"4D",x"2B",x"04",x"6E",x"9F",x"20",x"64",x"D6",x"E3",x"27",x"08",x"8D",x"D0",x"D3",x"7A",
    x"DD",x"7A",x"0F",x"E3",x"D6",x"E4",x"27",x"08",x"8D",x"C4",x"D3",x"7C",x"DD",x"7C",x"0F",x"E4",
    x"0C",x"31",x"96",x"31",x"84",x"03",x"26",x"41",x"0D",x"7E",x"27",x"0A",x"0A",x"7E",x"26",x"06",
    x"A6",x"C4",x"84",x"FB",x"A7",x"C4",x"D6",x"19",x"C5",x"04",x"27",x"1D",x"A6",x"C4",x"34",x"02",
    x"8A",x"01",x"A7",x"C4",x"96",x"77",x"2A",x"07",x"96",x"1C",x"44",x"25",x"02",x"6A",x"C4",x"63",
    x"9F",x"20",x"21",x"03",x"30",x"35",x"02",x"A7",x"C4",x"0D",x"37",x"27",x"0C",x"96",x"38",x"91",
    x"76",x"27",x"02",x"0C",x"38",x"C4",x"FD",x"D7",x"19",x"A6",x"41",x"0D",x"63",x"27",x"04",x"6E",
    x"9F",x"20",x"61",x"3B",x"2A",x"10",x"A6",x"4C",x"85",x"04",x"26",x"03",x"0C",x"E3",x"8C",x"0A",
    x"E3",x"A6",x"4E",x"48",x"2A",x"0F",x"A6",x"4C",x"85",x"08",x"26",x"03",x"0C",x"E4",x"8C",x"0A",
    x"E4",x"A6",x"4E",x"2B",x"E1",x"0D",x"7E",x"26",x"16",x"A6",x"4F",x"84",x"FB",x"A7",x"4F",x"E6",
    x"4D",x"8A",x"04",x"A7",x"4F",x"C5",x"04",x"26",x"0A",x"A6",x"C4",x"8A",x"04",x"A7",x"C4",x"86",
    x"05",x"97",x"7E",x"3B",x"B6",x"A7",x"E9",x"85",x"08",x"27",x"08",x"B6",x"A7",x"EA",x"84",x"F7",
    x"B7",x"A7",x"EA",x"3B",x"7F",x"22",x"00",x"B6",x"A7",x"C0",x"8A",x"20",x"B7",x"A7",x"C0",x"C1",
    x"04",x"26",x"07",x"86",x"04",x"B7",x"A7",x"CB",x"20",x"0C",x"C1",x"01",x"25",x"05",x"22",x"06",
    x"86",x"36",x"8C",x"86",x"06",x"8C",x"86",x"26",x"B7",x"A7",x"DD",x"86",x"06",x"97",x"86",x"6E",
    x"9F",x"EF",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"10",x"10",
    x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"50",x"28",x"14",x"00",x"28",x"28",x"FE",x"28",x"FE",
    x"28",x"28",x"00",x"10",x"FC",x"12",x"7C",x"90",x"7C",x"10",x"00",x"00",x"46",x"26",x"10",x"08",
    x"64",x"62",x"00",x"00",x"3A",x"4C",x"4A",x"30",x"48",x"30",x"00",x"00",x"00",x"00",x"00",x"18",
    x"0C",x"0C",x"00",x"00",x"08",x"10",x"10",x"10",x"10",x"08",x"00",x"00",x"10",x"08",x"08",x"08",
    x"08",x"10",x"00",x"00",x"54",x"38",x"6C",x"38",x"54",x"00",x"00",x"00",x"10",x"10",x"7C",x"10",
    x"10",x"00",x"00",x"00",x"10",x"0C",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"00",
    x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"20",x"10",x"08",
    x"04",x"02",x"01",x"00",x"3C",x"62",x"52",x"4A",x"46",x"3C",x"00",x"00",x"3C",x"08",x"08",x"28",
    x"18",x"08",x"00",x"00",x"7E",x"40",x"3C",x"02",x"42",x"3C",x"00",x"00",x"3C",x"42",x"02",x"1C",
    x"42",x"3C",x"00",x"00",x"04",x"7E",x"24",x"14",x"0C",x"04",x"00",x"00",x"3C",x"42",x"02",x"7C",
    x"40",x"7E",x"00",x"00",x"3C",x"42",x"42",x"7C",x"20",x"1C",x"00",x"00",x"40",x"20",x"10",x"08",
    x"04",x"7E",x"00",x"00",x"3C",x"42",x"42",x"3C",x"42",x"3C",x"00",x"00",x"38",x"04",x"3E",x"42",
    x"42",x"3C",x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"00",x"00",x"10",x"0C",x"00",x"0C",x"0C",
    x"00",x"00",x"00",x"00",x"08",x"10",x"20",x"20",x"10",x"08",x"00",x"00",x"00",x"7E",x"00",x"7E",
    x"00",x"00",x"00",x"00",x"10",x"08",x"04",x"04",x"08",x"10",x"00",x"00",x"08",x"00",x"08",x"04",
    x"22",x"1C",x"00",x"00",x"3E",x"5C",x"52",x"5E",x"42",x"3C",x"00",x"00",x"42",x"42",x"7E",x"42",
    x"24",x"18",x"00",x"00",x"7E",x"22",x"22",x"3C",x"22",x"7C",x"00",x"00",x"3C",x"42",x"40",x"40",
    x"42",x"3C",x"00",x"00",x"7C",x"22",x"22",x"22",x"22",x"7C",x"00",x"00",x"7E",x"40",x"40",x"78",
    x"40",x"7E",x"00",x"00",x"40",x"40",x"40",x"78",x"40",x"7E",x"00",x"00",x"3C",x"42",x"4E",x"40",
    x"42",x"3C",x"00",x"00",x"42",x"42",x"42",x"7E",x"42",x"42",x"00",x"00",x"38",x"10",x"10",x"10",
    x"10",x"38",x"00",x"00",x"3C",x"42",x"02",x"02",x"02",x"02",x"00",x"00",x"44",x"48",x"50",x"70",
    x"48",x"44",x"00",x"00",x"7E",x"40",x"40",x"40",x"40",x"40",x"00",x"00",x"42",x"42",x"42",x"5A",
    x"66",x"42",x"00",x"00",x"42",x"46",x"4A",x"52",x"62",x"42",x"00",x"00",x"3C",x"42",x"42",x"42",
    x"42",x"3C",x"00",x"00",x"40",x"40",x"7C",x"42",x"42",x"7C",x"00",x"00",x"3A",x"44",x"4A",x"42",
    x"42",x"3C",x"00",x"00",x"42",x"44",x"7C",x"42",x"42",x"7C",x"00",x"00",x"3C",x"42",x"02",x"3C",
    x"40",x"3C",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"7C",x"00",x"00",x"3C",x"42",x"42",x"42",
    x"42",x"42",x"00",x"00",x"18",x"24",x"24",x"42",x"42",x"42",x"00",x"00",x"42",x"66",x"5A",x"42",
    x"42",x"42",x"00",x"00",x"42",x"24",x"18",x"18",x"24",x"42",x"00",x"00",x"10",x"10",x"10",x"10",
    x"28",x"44",x"00",x"00",x"7E",x"20",x"10",x"08",x"04",x"7E",x"00",x"00",x"38",x"20",x"20",x"20",
    x"20",x"38",x"00",x"01",x"02",x"04",x"08",x"10",x"20",x"40",x"80",x"00",x"1C",x"04",x"04",x"04",
    x"04",x"1C",x"00",x"00",x"10",x"10",x"10",x"7C",x"38",x"10",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"3A",x"44",x"38",x"04",
    x"38",x"00",x"00",x"00",x"5C",x"62",x"42",x"62",x"5C",x"40",x"00",x"00",x"3C",x"42",x"40",x"42",
    x"3C",x"00",x"00",x"00",x"3A",x"46",x"42",x"46",x"3A",x"02",x"00",x"00",x"3C",x"40",x"7E",x"42",
    x"3C",x"00",x"00",x"00",x"10",x"10",x"7C",x"10",x"12",x"0C",x"00",x"3C",x"02",x"3A",x"46",x"46",
    x"3C",x"00",x"00",x"00",x"42",x"42",x"42",x"62",x"5C",x"40",x"00",x"00",x"1C",x"08",x"08",x"08",
    x"18",x"00",x"08",x"38",x"44",x"04",x"04",x"04",x"04",x"00",x"04",x"00",x"22",x"34",x"28",x"24",
    x"22",x"20",x"00",x"00",x"1C",x"08",x"08",x"08",x"08",x"18",x"00",x"00",x"92",x"92",x"92",x"DA",
    x"A4",x"00",x"00",x"00",x"22",x"22",x"22",x"32",x"4C",x"00",x"00",x"00",x"3C",x"42",x"42",x"42",
    x"3C",x"00",x"00",x"40",x"5C",x"62",x"42",x"62",x"5C",x"00",x"00",x"02",x"3A",x"46",x"46",x"46",
    x"3A",x"00",x"00",x"00",x"40",x"40",x"40",x"62",x"5C",x"00",x"00",x"00",x"7C",x"02",x"3C",x"40",
    x"3C",x"00",x"00",x"00",x"0C",x"12",x"10",x"10",x"38",x"10",x"00",x"00",x"3A",x"46",x"42",x"42",
    x"42",x"00",x"00",x"00",x"18",x"24",x"42",x"42",x"42",x"00",x"00",x"00",x"24",x"5A",x"42",x"42",
    x"42",x"00",x"00",x"00",x"42",x"24",x"18",x"24",x"42",x"00",x"00",x"3C",x"42",x"1A",x"66",x"42",
    x"42",x"00",x"00",x"00",x"7E",x"20",x"18",x"04",x"7E",x"00",x"00",x"0C",x"08",x"08",x"10",x"08",
    x"08",x"0C",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"30",x"10",x"10",x"08",x"10",
    x"10",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"70",x"50",x"70",x"00",x"18",x"3C",x"42",x"40",x"42",
    x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"30",x"00",x"00",x"00",x"00",x"00",
    x"00",x"18",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"18",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"66",x"34",x"08",x"C6",x"20",x"1F",x"9B",x"D6",x"19",x"34",x"04",x"CA",x"10",x"D7",
    x"19",x"0F",x"35",x"0F",x"29",x"7E",x"E9",x"00",x"96",x"5C",x"81",x"30",x"25",x"05",x"D6",x"5C",
    x"7E",x"F6",x"1E",x"0D",x"5D",x"26",x"46",x"3F",x"0C",x"34",x"06",x"8E",x"02",x"71",x"30",x"1F",
    x"26",x"FC",x"3F",x"0C",x"10",x"A3",x"E1",x"26",x"F0",x"C1",x"3A",x"27",x"36",x"D1",x"37",x"26",
    x"10",x"96",x"38",x"91",x"76",x"25",x"2E",x"86",x"02",x"95",x"19",x"26",x"28",x"BD",x"F8",x"DD",
    x"8C",x"0F",x"38",x"D7",x"37",x"C1",x"3A",x"25",x"01",x"5A",x"3F",x"08",x"04",x"44",x"24",x"18",
    x"C1",x"3A",x"25",x"05",x"8E",x"F6",x"88",x"E6",x"85",x"CA",x"80",x"20",x"27",x"D6",x"5D",x"4F",
    x"7E",x"F6",x"1C",x"0F",x"37",x"5F",x"20",x"79",x"C1",x"3F",x"26",x"0E",x"86",x"10",x"A8",x"C4",
    x"A7",x"C4",x"96",x"19",x"88",x"80",x"97",x"19",x"20",x"EB",x"9E",x"6D",x"E6",x"85",x"04",x"44",
    x"24",x"04",x"C4",x"BF",x"20",x"38",x"04",x"44",x"24",x"59",x"C1",x"05",x"26",x"04",x"C6",x"25",
    x"20",x"2C",x"C1",x"1D",x"25",x"28",x"C1",x"2F",x"22",x"0E",x"10",x"8E",x"F6",x"8F",x"E6",x"A5",
    x"C1",x"06",x"26",x"1A",x"C6",x"30",x"20",x"35",x"C1",x"39",x"22",x"08",x"A6",x"C4",x"85",x"10",
    x"27",x"0C",x"20",x"4D",x"C1",x"3F",x"22",x"08",x"10",x"8E",x"F6",x"83",x"E6",x"A5",x"20",x"5E",
    x"C1",x"5B",x"27",x"04",x"C1",x"5D",x"26",x"04",x"CB",x"20",x"20",x"52",x"C1",x"5E",x"27",x"07",
    x"5D",x"2A",x"4B",x"CB",x"05",x"20",x"47",x"C6",x"48",x"0D",x"5C",x"26",x"41",x"D7",x"5C",x"C6",
    x"16",x"20",x"3D",x"C1",x"05",x"27",x"28",x"A6",x"C4",x"85",x"10",x"26",x"1E",x"C1",x"41",x"25",
    x"08",x"C1",x"5A",x"22",x"16",x"CB",x"20",x"20",x"25",x"C1",x"30",x"25",x"0E",x"C1",x"39",x"22",
    x"1D",x"10",x"8E",x"F6",x"A2",x"C0",x"30",x"E6",x"A5",x"20",x"04",x"0D",x"5C",x"27",x"25",x"86",
    x"07",x"4A",x"27",x"0F",x"30",x"1D",x"E1",x"84",x"26",x"F7",x"EC",x"01",x"97",x"5D",x"0F",x"5C",
    x"E7",x"64",x"39",x"86",x"06",x"4A",x"27",x"F6",x"30",x"1D",x"E1",x"84",x"26",x"F7",x"EC",x"01",
    x"DD",x"5C",x"20",x"AB",x"C1",x"16",x"26",x"E6",x"0C",x"5C",x"20",x"E4",x"04",x"41",x"61",x"01",
    x"42",x"65",x"02",x"41",x"65",x"05",x"41",x"75",x"03",x"4B",x"63",x"00",x"00",x"30",x"00",x"00",
    x"4B",x"00",x"00",x"41",x"00",x"00",x"42",x"5E",x"00",x"43",x"00",x"00",x"48",x"00",x"00",x"02",
    x"16",x"00",x"0D",x"1E",x"43",x"0B",x"57",x"31",x"3D",x"41",x"24",x"51",x"56",x"08",x"58",x"32",
    x"2D",x"5A",x"3A",x"53",x"42",x"0A",x"20",x"33",x"30",x"45",x"50",x"44",x"4D",x"09",x"23",x"34",
    x"39",x"52",x"4F",x"46",x"4C",x"3E",x"3B",x"35",x"38",x"54",x"49",x"47",x"4B",x"1C",x"2C",x"36",
    x"37",x"59",x"55",x"48",x"4A",x"1D",x"4E",x"05",x"5E",x"29",x"5D",x"5B",x"00",x"C1",x"C2",x"C3",
    x"C4",x"C5",x"04",x"2A",x"01",x"22",x"27",x"28",x"5F",x"02",x"21",x"03",x"7F",x"0C",x"00",x"00",
    x"00",x"00",x"40",x"26",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"3F",x"5C",x"2F",x"2E",x"00",
    x"2B",x"3C",x"30",x"03",x"19",x"38",x"06",x"1A",x"D0",x"BD",x"FC",x"00",x"0D",x"77",x"2A",x"08",
    x"96",x"1C",x"44",x"25",x"03",x"7A",x"A7",x"C0",x"8E",x"FE",x"16",x"96",x"59",x"AD",x"96",x"0F",
    x"2F",x"0F",x"2E",x"39",x"C1",x"20",x"24",x"33",x"C1",x"07",x"25",x"F7",x"4F",x"58",x"8E",x"FE",
    x"10",x"6E",x"95",x"0F",x"59",x"C1",x"4B",x"27",x"16",x"C1",x"30",x"27",x"17",x"86",x"02",x"97",
    x"5B",x"86",x"05",x"9E",x"6D",x"30",x"1D",x"E1",x"02",x"27",x"0A",x"4A",x"26",x"F7",x"8C",x"86",
    x"80",x"97",x"5B",x"39",x"4F",x"1F",x"89",x"CA",x"80",x"20",x"39",x"96",x"77",x"27",x"15",x"2B",
    x"0B",x"BD",x"F8",x"EC",x"96",x"77",x"85",x"02",x"26",x"07",x"20",x"08",x"96",x"1C",x"44",x"25",
    x"03",x"BD",x"FC",x"09",x"0F",x"2F",x"0D",x"5B",x"2B",x"11",x"27",x"06",x"C1",x"61",x"24",x"14",
    x"0F",x"5B",x"5D",x"2A",x"0F",x"DE",x"70",x"C0",x"80",x"20",x"0D",x"C1",x"63",x"26",x"F1",x"D6",
    x"5B",x"5C",x"0F",x"5B",x"DE",x"73",x"C0",x"20",x"86",x"08",x"3D",x"33",x"CB",x"0F",x"30",x"10",
    x"9E",x"21",x"96",x"77",x"44",x"25",x"08",x"8E",x"F7",x"9C",x"CC",x"F7",x"B4",x"20",x"06",x"8E",
    x"F7",x"F0",x"CC",x"F7",x"C3",x"34",x"16",x"D6",x"2A",x"C4",x"03",x"54",x"10",x"26",x"00",x"BE",
    x"BD",x"F8",x"73",x"37",x"02",x"AD",x"F4",x"24",x"02",x"AD",x"F4",x"5A",x"26",x"F5",x"32",x"64",
    x"BD",x"F8",x"A7",x"8D",x"1F",x"30",x"1F",x"26",x"FA",x"7E",x"F8",x"6E",x"0D",x"77",x"2A",x"12",
    x"34",x"03",x"8D",x"16",x"44",x"25",x"03",x"E7",x"A4",x"8C",x"E7",x"21",x"8D",x"0C",x"35",x"03",
    x"20",x"02",x"E7",x"21",x"A7",x"A4",x"31",x"A8",x"D8",x"39",x"B6",x"A7",x"C0",x"88",x"01",x"B7",
    x"A7",x"C0",x"39",x"34",x"07",x"8E",x"F7",x"FE",x"96",x"2B",x"D6",x"2B",x"84",x"03",x"48",x"48",
    x"C4",x"30",x"3A",x"30",x"86",x"A6",x"61",x"A4",x"02",x"A8",x"03",x"A7",x"A4",x"7A",x"A7",x"C0",
    x"A6",x"61",x"A4",x"84",x"A8",x"01",x"A7",x"A4",x"7C",x"A7",x"C0",x"31",x"A8",x"D8",x"35",x"87",
    x"8D",x"D1",x"31",x"A8",x"29",x"1E",x"98",x"8D",x"CA",x"31",x"3F",x"1E",x"89",x"39",x"00",x"00",
    x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
    x"00",x"00",x"00",x"FF",x"00",x"00",x"FF",x"00",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"00",x"00",
    x"FF",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",
    x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"00",x"FF",x"00",x"FF",x"8D",x"33",
    x"37",x"02",x"34",x"05",x"97",x"44",x"CC",x"80",x"00",x"04",x"44",x"46",x"56",x"47",x"56",x"24",
    x"F8",x"35",x"01",x"AD",x"F8",x"03",x"24",x"03",x"AD",x"F8",x"03",x"35",x"04",x"5A",x"26",x"E0",
    x"32",x"64",x"8D",x"43",x"BD",x"F7",x"9C",x"30",x"1F",x"26",x"F9",x"8C",x"32",x"62",x"0D",x"5B",
    x"27",x"4D",x"39",x"C6",x"08",x"0D",x"5B",x"27",x"06",x"0A",x"5B",x"26",x"02",x"5A",x"5A",x"39",
    x"DE",x"2B",x"9E",x"21",x"10",x"9E",x"1B",x"96",x"2A",x"C6",x"FF",x"D7",x"2C",x"C6",x"20",x"3F",
    x"02",x"D6",x"1C",x"C1",x"01",x"26",x"F6",x"DF",x"2B",x"9F",x"21",x"10",x"9F",x"1B",x"97",x"2A",
    x"86",x"FF",x"A7",x"9F",x"20",x"1A",x"39",x"8E",x"00",x"08",x"24",x"02",x"30",x"08",x"86",x"40",
    x"94",x"19",x"26",x"B8",x"10",x"9E",x"21",x"BD",x"FC",x"09",x"96",x"2B",x"D6",x"2B",x"39",x"96",
    x"2A",x"85",x"02",x"27",x"04",x"0C",x"1C",x"0C",x"22",x"20",x"67",x"8D",x"1F",x"86",x"FB",x"20",
    x"06",x"0D",x"77",x"26",x"0C",x"86",x"BF",x"94",x"19",x"20",x"04",x"86",x"40",x"9A",x"19",x"97",
    x"19",x"39",x"A6",x"64",x"84",x"EF",x"A7",x"64",x"86",x"04",x"20",x"F1",x"96",x"19",x"85",x"04",
    x"27",x"19",x"0D",x"30",x"27",x"15",x"BD",x"FC",x"00",x"0D",x"77",x"2A",x"08",x"96",x"1C",x"44",
    x"25",x"03",x"7A",x"A7",x"C0",x"63",x"9F",x"20",x"21",x"03",x"30",x"39",x"8D",x"DE",x"0F",x"1C",
    x"0C",x"1C",x"BD",x"F9",x"98",x"20",x"89",x"8D",x"D3",x"0C",x"1B",x"96",x"1B",x"91",x"20",x"23",
    x"77",x"5F",x"20",x"59",x"8D",x"C6",x"0F",x"1C",x"0C",x"1C",x"20",x"68",x"8D",x"28",x"86",x"FF",
    x"97",x"2E",x"0C",x"1C",x"96",x"1C",x"0D",x"77",x"2B",x"0A",x"81",x"29",x"27",x"21",x"81",x"2A",
    x"27",x"1B",x"20",x"08",x"81",x"51",x"27",x"17",x"81",x"52",x"27",x"11",x"0D",x"2F",x"27",x"03",
    x"BD",x"F9",x"D9",x"7E",x"FD",x"76",x"8D",x"94",x"9E",x"21",x"C6",x"08",x"39",x"0A",x"22",x"0D",
    x"2F",x"27",x"07",x"31",x"89",x"01",x"19",x"BD",x"F9",x"ED",x"CC",x"01",x"01",x"97",x"1C",x"0D",
    x"2E",x"2B",x"0A",x"9E",x"1A",x"D5",x"2A",x"27",x"02",x"6F",x"1F",x"6F",x"84",x"D4",x"2A",x"58",
    x"58",x"58",x"8E",x"FE",x"50",x"3A",x"96",x"1B",x"AB",x"84",x"97",x"1B",x"91",x"20",x"23",x"08",
    x"0D",x"2C",x"27",x"07",x"96",x"1E",x"97",x"1B",x"7E",x"FD",x"76",x"9F",x"44",x"E6",x"84",x"10",
    x"9E",x"1D",x"10",x"9C",x"1F",x"24",x"06",x"A6",x"21",x"A7",x"A0",x"20",x"F5",x"86",x"FF",x"A7",
    x"A4",x"5A",x"26",x"EB",x"A6",x"84",x"48",x"48",x"48",x"8E",x"FA",x"FC",x"CE",x"FB",x"1F",x"BD",
    x"FA",x"70",x"20",x"7A",x"0D",x"77",x"2A",x"0D",x"BD",x"FC",x"00",x"96",x"1C",x"44",x"25",x"05",
    x"7A",x"A7",x"C0",x"20",x"16",x"31",x"1F",x"20",x"14",x"0D",x"77",x"2A",x"0B",x"BD",x"FC",x"00",
    x"96",x"1C",x"44",x"24",x"06",x"7A",x"A7",x"C0",x"31",x"01",x"8C",x"31",x"84",x"A6",x"84",x"8D",
    x"0C",x"30",x"88",x"D8",x"BD",x"F7",x"B4",x"8D",x"04",x"5A",x"26",x"F1",x"39",x"34",x"02",x"0D",
    x"77",x"2A",x"03",x"BD",x"F7",x"BA",x"35",x"82",x"BD",x"F9",x"56",x"96",x"1C",x"81",x"01",x"2E",
    x"17",x"0D",x"2F",x"27",x"06",x"31",x"89",x"FE",x"E7",x"8D",x"D2",x"C6",x"28",x"0D",x"77",x"2A",
    x"01",x"58",x"D7",x"1C",x"8D",x"0A",x"20",x"0E",x"0D",x"2F",x"27",x"02",x"8D",x"96",x"0A",x"1C",
    x"7E",x"FD",x"76",x"BD",x"F8",x"EC",x"96",x"1B",x"91",x"1E",x"2F",x"07",x"4A",x"8C",x"96",x"20",
    x"7E",x"F9",x"96",x"0D",x"2C",x"26",x"F7",x"CC",x"08",x"01",x"D4",x"2A",x"27",x"01",x"48",x"34",
    x"02",x"10",x"9E",x"1F",x"10",x"9C",x"1D",x"23",x"06",x"E6",x"A2",x"E7",x"21",x"20",x"F5",x"C6",
    x"FF",x"E7",x"A4",x"44",x"85",x"08",x"26",x"E9",x"35",x"02",x"8E",x"FA",x"B2",x"CE",x"FA",x"DD",
    x"34",x"52",x"6A",x"E4",x"2B",x"3A",x"BD",x"FC",x"00",x"96",x"77",x"85",x"02",x"27",x"03",x"7A",
    x"A7",x"C0",x"AD",x"F8",x"01",x"DC",x"27",x"AD",x"F8",x"03",x"96",x"2B",x"34",x"02",x"96",x"77",
    x"85",x"C1",x"26",x"07",x"86",x"40",x"94",x"19",x"26",x"0E",x"8C",x"0F",x"2B",x"3F",x"04",x"AD",
    x"F8",x"02",x"BD",x"F8",x"BA",x"AD",x"F8",x"04",x"35",x"02",x"97",x"2B",x"0D",x"2D",x"26",x"C2",
    x"35",x"D2",x"10",x"DF",x"46",x"DC",x"23",x"C3",x"00",x"28",x"DD",x"44",x"DE",x"25",x"32",x"C8",
    x"D1",x"0D",x"2D",x"26",x"04",x"32",x"E9",x"FE",x"E8",x"35",x"3E",x"36",x"3E",x"32",x"72",x"11",
    x"B3",x"20",x"44",x"22",x"F4",x"86",x"20",x"1F",x"8B",x"10",x"DE",x"46",x"39",x"10",x"DF",x"46",
    x"1F",x"01",x"1F",x"02",x"1F",x"04",x"DE",x"23",x"33",x"C8",x"28",x"0D",x"2D",x"26",x"04",x"33",
    x"C9",x"01",x"18",x"36",x"76",x"11",x"93",x"23",x"22",x"F9",x"20",x"DD",x"10",x"DF",x"46",x"10",
    x"DE",x"44",x"EC",x"65",x"DE",x"23",x"32",x"C8",x"28",x"33",x"47",x"0D",x"2D",x"26",x"02",x"32",
    x"EB",x"35",x"3E",x"36",x"3E",x"33",x"4E",x"11",x"BC",x"20",x"25",x"25",x"F4",x"20",x"B6",x"10",
    x"DF",x"46",x"1F",x"01",x"1F",x"02",x"10",x"DE",x"44",x"EC",x"63",x"DE",x"25",x"33",x"C8",x"E0",
    x"0D",x"2D",x"26",x"02",x"33",x"CB",x"1F",x"10",x"1F",x"04",x"36",x"76",x"33",x"C8",x"10",x"11",
    x"93",x"25",x"23",x"F6",x"20",x"93",x"BD",x"FC",x"00",x"96",x"77",x"85",x"02",x"27",x"03",x"7A",
    x"A7",x"C0",x"0F",x"30",x"D6",x"2B",x"34",x"04",x"DC",x"27",x"1F",x"01",x"1F",x"02",x"DE",x"25",
    x"36",x"36",x"36",x"30",x"11",x"93",x"23",x"2E",x"F7",x"96",x"77",x"85",x"E1",x"26",x"07",x"86",
    x"40",x"94",x"19",x"26",x"0F",x"8C",x"0F",x"2B",x"C6",x"01",x"F4",x"A7",x"C0",x"27",x"05",x"BD",
    x"F8",x"B7",x"20",x"D6",x"35",x"04",x"D7",x"2B",x"9E",x"1D",x"86",x"FF",x"A7",x"80",x"9C",x"1F",
    x"23",x"FA",x"7E",x"F9",x"26",x"A6",x"64",x"1F",x"8A",x"96",x"19",x"85",x"08",x"26",x"0D",x"4F",
    x"B7",x"A7",x"C1",x"4C",x"5F",x"5C",x"2A",x"FD",x"81",x"11",x"26",x"F4",x"39",x"B6",x"A7",x"C3",
    x"84",x"F7",x"20",x"05",x"B6",x"A7",x"C3",x"8A",x"08",x"B7",x"A7",x"C3",x"39",x"C4",x"03",x"96",
    x"2A",x"84",x"FC",x"8D",x"2B",x"97",x"2A",x"39",x"0D",x"77",x"26",x"28",x"9E",x"23",x"3F",x"04",
    x"A6",x"84",x"8D",x"14",x"A7",x"80",x"9C",x"25",x"26",x"F6",x"96",x"77",x"27",x"03",x"44",x"24",
    x"13",x"96",x"2B",x"8D",x"03",x"7E",x"FC",x"6B",x"1F",x"89",x"44",x"44",x"44",x"44",x"8D",x"27",
    x"34",x"04",x"AB",x"E0",x"39",x"C4",x"0F",x"D7",x"86",x"FA",x"A7",x"E4",x"F7",x"A7",x"DD",x"39",
    x"34",x"02",x"86",x"01",x"BA",x"A7",x"C0",x"20",x"07",x"34",x"02",x"86",x"FE",x"B4",x"A7",x"C0",
    x"B7",x"A7",x"C0",x"35",x"82",x"86",x"0F",x"58",x"58",x"58",x"58",x"39",x"0D",x"77",x"26",x"2F",
    x"C4",x"0F",x"86",x"F0",x"34",x"02",x"8D",x"0F",x"35",x"02",x"C4",x"0F",x"96",x"77",x"27",x"03",
    x"44",x"24",x"1C",x"86",x"F0",x"20",x"30",x"3F",x"04",x"D7",x"44",x"D7",x"45",x"9E",x"23",x"EC",
    x"84",x"A4",x"62",x"E4",x"62",x"D3",x"44",x"ED",x"81",x"9C",x"25",x"26",x"F2",x"D6",x"44",x"39",
    x"0D",x"77",x"26",x"FB",x"8D",x"BF",x"34",x"02",x"8D",x"DD",x"35",x"02",x"20",x"09",x"96",x"77",
    x"27",x"03",x"44",x"24",x"EA",x"8D",x"AE",x"94",x"2B",x"8D",x"85",x"97",x"2B",x"39",x"0F",x"2C",
    x"C1",x"7A",x"27",x"08",x"0F",x"2D",x"54",x"24",x"05",x"03",x"2D",x"8C",x"03",x"2C",x"39",x"4C",
    x"4C",x"4C",x"48",x"97",x"59",x"39",x"96",x"77",x"27",x"1F",x"0F",x"77",x"5F",x"86",x"AF",x"94",
    x"19",x"97",x"19",x"F7",x"A7",x"DC",x"CC",x"00",x"00",x"DD",x"23",x"CC",x"1F",x"40",x"DD",x"25",
    x"0F",x"1E",x"86",x"18",x"97",x"20",x"BD",x"FB",x"46",x"39",x"C6",x"80",x"D5",x"77",x"26",x"F9",
    x"D7",x"77",x"C6",x"2A",x"86",x"50",x"9A",x"19",x"20",x"D7",x"C6",x"01",x"D5",x"77",x"26",x"E9",
    x"D7",x"77",x"C6",x"21",x"20",x"EE",x"C6",x"40",x"D5",x"77",x"26",x"DD",x"D7",x"77",x"C6",x"7B",
    x"20",x"E2",x"96",x"77",x"34",x"02",x"1F",x"98",x"44",x"25",x"03",x"86",x"02",x"8C",x"86",x"04",
    x"C0",x"82",x"2B",x"03",x"8B",x"08",x"5F",x"97",x"77",x"34",x"04",x"C6",x"26",x"EB",x"E0",x"86",
    x"0E",x"A4",x"E0",x"27",x"04",x"F7",x"A7",x"DC",x"39",x"96",x"77",x"34",x"02",x"86",x"80",x"97",
    x"77",x"8D",x"B1",x"35",x"02",x"97",x"77",x"39",x"C4",x"03",x"96",x"79",x"84",x"FC",x"34",x"04",
    x"AB",x"E0",x"97",x"79",x"C6",x"20",x"D5",x"77",x"26",x"8F",x"D7",x"77",x"C6",x"3F",x"20",x"D9",
    x"0D",x"5A",x"26",x"03",x"D7",x"5A",x"39",x"BD",x"F8",x"EC",x"C1",x"40",x"25",x"17",x"0D",x"77",
    x"2A",x"05",x"C8",x"C0",x"C4",x"7F",x"8C",x"C4",x"3F",x"D7",x"1C",x"D6",x"5A",x"C4",x"3F",x"D7",
    x"1B",x"8D",x"33",x"20",x"2C",x"C1",x"30",x"2C",x"28",x"DE",x"1B",x"9E",x"21",x"34",x"50",x"C1",
    x"20",x"2D",x"0D",x"8D",x"44",x"D7",x"1E",x"8D",x"1D",x"83",x"01",x"18",x"DD",x"23",x"20",x"0B",
    x"8D",x"37",x"D7",x"20",x"8D",x"10",x"C3",x"00",x"28",x"DD",x"25",x"35",x"50",x"DF",x"1B",x"9F",
    x"21",x"0F",x"5A",x"0F",x"59",x"39",x"96",x"1B",x"BD",x"FF",x"15",x"DD",x"21",x"0D",x"77",x"2A",
    x"12",x"BD",x"FC",x"09",x"D6",x"1C",x"54",x"24",x"04",x"7C",x"A7",x"C0",x"5C",x"4F",x"D3",x"21",
    x"DD",x"21",x"39",x"96",x"21",x"DB",x"1C",x"20",x"F7",x"0F",x"1C",x"0C",x"1C",x"C4",x"0F",x"D7",
    x"1B",x"96",x"5A",x"84",x"0F",x"C6",x"0A",x"3D",x"DB",x"1B",x"D7",x"1B",x"39",x"86",x"80",x"C1",
    x"20",x"27",x"1C",x"C1",x"40",x"25",x"1C",x"CE",x"FD",x"D4",x"0D",x"2A",x"2B",x"02",x"33",x"4F",
    x"E1",x"C4",x"33",x"43",x"25",x"FA",x"AD",x"D3",x"0F",x"59",x"86",x"7F",x"94",x"2A",x"8C",x"9A",
    x"2A",x"97",x"2A",x"39",x"7C",x"FD",x"C8",x"7B",x"FB",x"C8",x"60",x"FD",x"C8",x"50",x"FC",x"1C",
    x"40",x"FC",x"50",x"88",x"FD",x"C8",x"84",x"FD",x"08",x"80",x"FC",x"D2",x"7F",x"FC",x"C6",x"7E",
    x"FC",x"BA",x"7D",x"FC",x"AA",x"7C",x"FC",x"86",x"7B",x"FB",x"DA",x"78",x"FC",x"6E",x"77",x"FB",
    x"AD",x"76",x"FB",x"B4",x"75",x"F8",x"DB",x"74",x"F8",x"D1",x"70",x"FB",x"BD",x"60",x"FB",x"F5",
    x"50",x"FC",x"2A",x"40",x"FC",x"5E",x"F6",x"E4",x"FD",x"AD",x"FD",x"20",x"F6",x"F3",x"FB",x"95",
    x"FA",x"08",x"F9",x"2C",x"F9",x"17",x"FA",x"33",x"FB",x"46",x"F9",x"0C",x"F6",x"E3",x"F6",x"E3",
    x"F6",x"E3",x"F8",x"E2",x"F6",x"E3",x"F6",x"E3",x"F8",x"CB",x"F6",x"E3",x"FC",x"7F",x"F6",x"E3",
    x"F8",x"80",x"F6",x"E3",x"F6",x"E3",x"FC",x"81",x"F6",x"E3",x"F6",x"E3",x"F9",x"24",x"FC",x"80",
    x"01",x"01",x"19",x"FE",x"E8",x"01",x"18",x"00",x"02",x"02",x"59",x"FD",x"A8",x"02",x"58",x"01",
    x"D6",x"19",x"34",x"04",x"C6",x"14",x"3F",x"02",x"0D",x"5D",x"10",x"2E",x"00",x"90",x"10",x"2B",
    x"00",x"94",x"C6",x"1F",x"E7",x"65",x"BD",x"FF",x"15",x"0D",x"77",x"27",x"23",x"1F",x"03",x"BD",
    x"FC",x"09",x"E6",x"68",x"96",x"77",x"85",x"80",x"27",x"0C",x"57",x"24",x"04",x"5C",x"7C",x"A7",
    x"C0",x"4F",x"33",x"CB",x"20",x"0E",x"85",x"0E",x"27",x"F4",x"85",x"04",x"27",x"F3",x"20",x"EE",
    x"EB",x"68",x"1F",x"03",x"9E",x"73",x"CC",x"62",x"08",x"8D",x"73",x"25",x"3B",x"30",x"06",x"33",
    x"C9",x"FF",x"10",x"64",x"65",x"CC",x"04",x"02",x"8D",x"64",x"24",x"4C",x"E6",x"65",x"C1",x"44",
    x"26",x"02",x"C6",x"48",x"D7",x"5D",x"C6",x"60",x"E7",x"65",x"9E",x"73",x"30",x"89",x"02",x"08",
    x"33",x"C9",x"00",x"F0",x"CC",x"1B",x"06",x"8D",x"45",x"25",x"03",x"C6",x"20",x"8C",x"E6",x"65",
    x"D7",x"5C",x"C6",x"16",x"E7",x"65",x"20",x"28",x"6D",x"65",x"2A",x"1E",x"C6",x"16",x"64",x"65",
    x"E7",x"65",x"25",x"05",x"CC",x"80",x"30",x"20",x"13",x"CC",x"4B",x"63",x"20",x"0E",x"D6",x"5D",
    x"E7",x"65",x"86",x"80",x"20",x"08",x"96",x"5C",x"A7",x"65",x"DC",x"27",x"D7",x"5C",x"97",x"5D",
    x"35",x"02",x"97",x"19",x"39",x"C6",x"A0",x"3D",x"58",x"49",x"C3",x"01",x"17",x"39",x"34",x"56",
    x"A6",x"80",x"A1",x"C4",x"26",x"08",x"33",x"C8",x"D8",x"5A",x"26",x"F4",x"43",x"21",x"4F",x"35",
    x"56",x"6C",x"67",x"30",x"08",x"25",x"03",x"4A",x"26",x"E4",x"39",x"43",x"53",x"C3",x"00",x"01",
    x"39",x"20",x"10",x"08",x"04",x"02",x"01",x"B6",x"A7",x"E4",x"BA",x"20",x"86",x"34",x"02",x"8A",
    x"30",x"B7",x"A7",x"DD",x"B6",x"A7",x"E6",x"85",x"20",x"27",x"22",x"34",x"02",x"7F",x"A7",x"E6",
    x"7F",x"A7",x"CB",x"A6",x"63",x"BD",x"B0",x"00",x"35",x"02",x"B7",x"A7",x"E6",x"44",x"44",x"44",
    x"B8",x"A7",x"E6",x"84",x"0C",x"B8",x"A7",x"E6",x"B7",x"A7",x"CB",x"20",x"05",x"A6",x"62",x"BD",
    x"B0",x"00",x"35",x"02",x"B7",x"A7",x"DD",x"E7",x"62",x"3B",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"35",x"40",x"DF",x"82",x"A6",
    x"C4",x"97",x"80",x"39",x"BD",x"CB",x"ED",x"8D",x"03",x"BD",x"CB",x"83",x"7E",x"CB",x"F9",x"FF",
    x"01",x"00",x"F0",x"53",x"FF",x"47",x"F0",x"A1",x"F0",x"B9",x"F0",x"9D",x"F0",x"53",x"F1",x"97");

  CONSTANT ROM_MO6_1 : arr8 := (
    x"A6",x"E4",x"84",x"F0",x"A7",x"E4",x"1F",x"8A",x"86",x"20",x"1F",x"8B",x"E6",x"F8",x"0A",x"C4",
    x"7F",x"CE",x"A7",x"C0",x"9E",x"6A",x"EC",x"85",x"85",x"F0",x"27",x"0F",x"8E",x"F0",x"37",x"8A",
    x"00",x"34",x"16",x"A6",x"C4",x"84",x"DF",x"A7",x"C4",x"20",x"07",x"8E",x"F0",x"43",x"8A",x"F0",
    x"34",x"16",x"EC",x"65",x"AE",x"68",x"39",x"34",x"01",x"B6",x"A7",x"C0",x"84",x"DF",x"B7",x"A7",
    x"C0",x"35",x"01",x"1F",x"A8",x"84",x"8F",x"AA",x"E4",x"A7",x"E4",x"AE",x"6A",x"E6",x"80",x"2B",
    x"03",x"AF",x"6A",x"3B",x"35",x"7F",x"32",x"62",x"39",x"01",x"9F",x"F6",x"C7",x"FC",x"09",x"FC",
    x"00",x"FB",x"99",x"F5",x"08",x"02",x"C3",x"06",x"69",x"04",x"A3",x"04",x"C1",x"04",x"E7",x"07",
    x"FA",x"08",x"24",x"FE",x"60",x"0A",x"C1",x"09",x"5A",x"03",x"44",x"04",x"64",x"09",x"D2",x"A0",
    x"04",x"A0",x"07",x"A0",x"0A",x"A0",x"1C",x"A0",x"19",x"A0",x"16",x"A0",x"22",x"A0",x"0D",x"A0",
    x"1F",x"A0",x"10",x"A0",x"13",x"0C",x"71",x"0C",x"E2",x"0C",x"F7",x"0A",x"E7",x"6E",x"9F",x"20",
    x"5E",x"6E",x"9F",x"20",x"67",x"3B",x"3B",x"3B",x"3B",x"3B",x"3B",x"3B",x"3B",x"3B",x"C1",x"05",
    x"23",x"05",x"C1",x"FB",x"24",x"01",x"58",x"1D",x"39",x"C6",x"20",x"1F",x"9B",x"CE",x"A7",x"C0",
    x"96",x"79",x"48",x"2A",x"06",x"A6",x"4E",x"85",x"C0",x"26",x"79",x"A6",x"43",x"85",x"01",x"27",
    x"03",x"4D",x"2B",x"04",x"6E",x"9F",x"20",x"64",x"D6",x"E3",x"27",x"08",x"8D",x"D0",x"D3",x"7A",
    x"DD",x"7A",x"0F",x"E3",x"D6",x"E4",x"27",x"08",x"8D",x"C4",x"D3",x"7C",x"DD",x"7C",x"0F",x"E4",
    x"0C",x"31",x"96",x"31",x"84",x"03",x"26",x"41",x"0D",x"7E",x"27",x"0A",x"0A",x"7E",x"26",x"06",
    x"A6",x"C4",x"84",x"FB",x"A7",x"C4",x"D6",x"19",x"C5",x"04",x"27",x"1D",x"A6",x"C4",x"34",x"02",
    x"8A",x"01",x"A7",x"C4",x"96",x"77",x"2A",x"07",x"96",x"1C",x"44",x"25",x"02",x"6A",x"C4",x"63",
    x"9F",x"20",x"21",x"03",x"30",x"35",x"02",x"A7",x"C4",x"0D",x"37",x"27",x"0C",x"96",x"38",x"91",
    x"76",x"27",x"02",x"0C",x"38",x"C4",x"FD",x"D7",x"19",x"A6",x"41",x"0D",x"63",x"27",x"04",x"6E",
    x"9F",x"20",x"61",x"3B",x"2A",x"10",x"A6",x"4C",x"85",x"04",x"26",x"03",x"0C",x"E3",x"8C",x"0A",
    x"E3",x"A6",x"4E",x"48",x"2A",x"0F",x"A6",x"4C",x"85",x"08",x"26",x"03",x"0C",x"E4",x"8C",x"0A",
    x"E4",x"A6",x"4E",x"2B",x"E1",x"0D",x"7E",x"26",x"16",x"A6",x"4F",x"84",x"FB",x"A7",x"4F",x"E6",
    x"4D",x"8A",x"04",x"A7",x"4F",x"C5",x"04",x"26",x"0A",x"A6",x"C4",x"8A",x"04",x"A7",x"C4",x"86",
    x"05",x"97",x"7E",x"3B",x"B6",x"A7",x"E9",x"85",x"08",x"27",x"08",x"B6",x"A7",x"EA",x"84",x"F7",
    x"B7",x"A7",x"EA",x"3B",x"47",x"75",x"79",x"B6",x"A7",x"C0",x"84",x"DF",x"B7",x"A7",x"C0",x"C6",
    x"20",x"1F",x"9B",x"10",x"CE",x"20",x"CC",x"CE",x"A5",x"5A",x"11",x"93",x"FE",x"27",x"1A",x"DF",
    x"FE",x"DF",x"7F",x"CC",x"07",x"0C",x"97",x"76",x"4F",x"DD",x"77",x"0F",x"79",x"8E",x"F2",x"93",
    x"86",x"FF",x"BD",x"FC",x"71",x"C6",x"20",x"1F",x"9B",x"B6",x"A7",x"DA",x"8E",x"A0",x"00",x"A6",
    x"84",x"81",x"52",x"26",x"06",x"96",x"80",x"81",x"5A",x"26",x"1E",x"0F",x"80",x"86",x"55",x"AB",
    x"80",x"AB",x"80",x"AB",x"80",x"A1",x"84",x"26",x"10",x"03",x"80",x"B6",x"A0",x"00",x"81",x"52",
    x"27",x"07",x"86",x"01",x"97",x"48",x"BD",x"A0",x"04",x"4F",x"8E",x"20",x"76",x"CE",x"F2",x"B3",
    x"37",x"20",x"A7",x"82",x"10",x"AF",x"83",x"8C",x"20",x"5E",x"2E",x"F4",x"A7",x"82",x"8C",x"20",
    x"19",x"2E",x"F9",x"43",x"A7",x"82",x"8C",x"20",x"00",x"2E",x"F9",x"D7",x"1A",x"D7",x"1D",x"D7",
    x"1F",x"CE",x"A7",x"C0",x"4F",x"5F",x"ED",x"42",x"ED",x"4E",x"ED",x"4C",x"86",x"7F",x"A7",x"41",
    x"86",x"04",x"A7",x"42",x"86",x"30",x"A7",x"C4",x"0F",x"7E",x"6F",x"42",x"86",x"75",x"A7",x"C4",
    x"8E",x"3E",x"3F",x"AF",x"42",x"8E",x"04",x"34",x"AF",x"4E",x"96",x"79",x"85",x"40",x"27",x"03",
    x"BD",x"FD",x"15",x"4F",x"B7",x"A7",x"E4",x"C6",x"26",x"FD",x"A7",x"DC",x"7F",x"A7",x"E6",x"86",
    x"93",x"B7",x"A7",x"E7",x"97",x"81",x"86",x"02",x"B7",x"A7",x"E5",x"86",x"04",x"9A",x"19",x"97",
    x"19",x"CC",x"1F",x"40",x"DD",x"25",x"86",x"18",x"97",x"20",x"B6",x"A0",x"00",x"81",x"52",x"26",
    x"0C",x"B6",x"22",x"8D",x"81",x"7E",x"26",x"05",x"C6",x"02",x"7E",x"F1",x"97",x"1C",x"EF",x"6E",
    x"9F",x"EF",x"FE",x"00",x"00",x"10",x"0F",x"10",x"F0",x"10",x"FF",x"1F",x"00",x"1F",x"0F",x"1F",
    x"F0",x"1F",x"FF",x"17",x"77",x"13",x"3A",x"13",x"A3",x"13",x"AA",x"1A",x"33",x"1A",x"3A",x"1E",
    x"E7",x"10",x"7B",x"F1",x"C3",x"F1",x"C3",x"F6",x"5D",x"F0",x"59",x"F0",x"53",x"F0",x"53",x"F0",
    x"53",x"F0",x"00",x"DC",x"27",x"DD",x"44",x"C6",x"72",x"E7",x"41",x"A6",x"41",x"2B",x"12",x"86",
    x"01",x"C1",x"72",x"27",x"0A",x"48",x"C1",x"6A",x"27",x"05",x"48",x"C1",x"70",x"26",x"58",x"97",
    x"44",x"0C",x"45",x"C0",x"02",x"2A",x"E2",x"0C",x"45",x"1F",x"A8",x"34",x"02",x"1A",x"50",x"A6",
    x"C4",x"84",x"F7",x"A7",x"C4",x"A6",x"42",x"34",x"02",x"84",x"FB",x"A7",x"42",x"A6",x"C4",x"8A",
    x"08",x"A7",x"C4",x"C6",x"40",x"E7",x"41",x"A6",x"41",x"2A",x"06",x"0C",x"45",x"C0",x"10",x"2A",
    x"F4",x"A6",x"C4",x"84",x"F7",x"A7",x"C4",x"35",x"02",x"8A",x"04",x"A7",x"42",x"35",x"02",x"1F",
    x"8A",x"D6",x"45",x"C1",x"40",x"26",x"10",x"C6",x"74",x"E7",x"41",x"A6",x"41",x"2A",x"08",x"0C",
    x"45",x"CB",x"02",x"C5",x"0E",x"26",x"F2",x"DC",x"44",x"C1",x"46",x"26",x"02",x"C6",x"3A",x"ED",
    x"63",x"C1",x"3A",x"39",x"1A",x"D0",x"6D",x"63",x"10",x"27",x"00",x"D3",x"A6",x"C4",x"97",x"44",
    x"A6",x"C4",x"98",x"44",x"2A",x"FA",x"03",x"44",x"C6",x"05",x"8E",x"00",x"00",x"A6",x"C4",x"98",
    x"44",x"2B",x"04",x"30",x"01",x"20",x"F6",x"03",x"44",x"34",x"10",x"5A",x"26",x"EC",x"C6",x"05",
    x"35",x"10",x"8C",x"00",x"10",x"25",x"2A",x"8C",x"00",x"1A",x"25",x"0C",x"8C",x"00",x"25",x"25",
    x"20",x"8C",x"00",x"33",x"25",x"07",x"20",x"19",x"8E",x"01",x"A1",x"20",x"03",x"8E",x"03",x"41",
    x"C1",x"05",x"27",x"06",x"9C",x"44",x"27",x"04",x"20",x"07",x"9F",x"44",x"5A",x"26",x"D1",x"20",
    x"07",x"5A",x"27",x"A8",x"35",x"10",x"20",x"F9",x"8C",x"01",x"A1",x"26",x"05",x"8E",x"00",x"24",
    x"20",x"03",x"8E",x"00",x"41",x"34",x"10",x"A6",x"C4",x"C6",x"FF",x"DD",x"44",x"32",x"7E",x"8D",
    x"3C",x"4D",x"26",x"FB",x"8D",x"37",x"96",x"45",x"81",x"01",x"26",x"F8",x"32",x"62",x"8D",x"45",
    x"81",x"01",x"27",x"FA",x"81",x"3C",x"27",x"05",x"32",x"62",x"7E",x"F3",x"4C",x"8D",x"36",x"81",
    x"5A",x"26",x"F5",x"8D",x"30",x"A7",x"66",x"8D",x"2C",x"A7",x"A0",x"97",x"41",x"6F",x"65",x"0A",
    x"41",x"27",x"6E",x"8D",x"20",x"A7",x"A0",x"AB",x"65",x"A7",x"65",x"20",x"F2",x"A6",x"C4",x"98",
    x"44",x"2A",x"FA",x"AE",x"64",x"8D",x"6E",x"A6",x"C4",x"98",x"44",x"2A",x"04",x"03",x"44",x"4F",
    x"21",x"43",x"09",x"45",x"39",x"C6",x"08",x"8D",x"E4",x"5A",x"26",x"FB",x"96",x"45",x"39",x"86",
    x"04",x"95",x"79",x"26",x"08",x"8E",x"00",x"13",x"CC",x"00",x"17",x"20",x"06",x"8E",x"00",x"2C",
    x"CC",x"00",x"32",x"34",x"16",x"CC",x"01",x"10",x"DD",x"40",x"96",x"40",x"8D",x"44",x"0A",x"41",
    x"26",x"F8",x"86",x"3C",x"8D",x"3C",x"86",x"5A",x"8D",x"38",x"A6",x"68",x"8D",x"34",x"A6",x"A4",
    x"97",x"41",x"A6",x"A0",x"8D",x"2C",x"0A",x"41",x"26",x"F8",x"32",x"62",x"8E",x"08",x"00",x"8D",
    x"14",x"32",x"62",x"39",x"E6",x"42",x"44",x"24",x"12",x"C4",x"F7",x"E7",x"42",x"44",x"24",x"0A",
    x"8D",x"00",x"8E",x"96",x"3D",x"30",x"1F",x"26",x"FC",x"4F",x"39",x"CA",x"08",x"8D",x"F3",x"E7",
    x"42",x"39",x"97",x"45",x"C6",x"08",x"8D",x"14",x"AE",x"64",x"8D",x"E9",x"AE",x"62",x"08",x"45",
    x"24",x"04",x"8D",x"08",x"30",x"1D",x"8D",x"DD",x"5A",x"26",x"EB",x"39",x"86",x"40",x"A8",x"C4",
    x"A7",x"C4",x"39",x"7D",x"20",x"36",x"26",x"19",x"34",x"7E",x"8D",x"0B",x"BD",x"F5",x"7E",x"BD",
    x"F5",x"46",x"BD",x"F6",x"07",x"35",x"FE",x"86",x"20",x"1F",x"8B",x"9F",x"32",x"10",x"9F",x"34",
    x"39",x"34",x"0E",x"8D",x"F2",x"96",x"2C",x"34",x"02",x"8A",x"80",x"97",x"2C",x"C6",x"1F",x"3F",
    x"02",x"1F",x"20",x"CB",x"40",x"3F",x"02",x"1F",x"10",x"CB",x"40",x"3F",x"02",x"D6",x"36",x"3F",
    x"02",x"35",x"02",x"97",x"2C",x"35",x"8E",x"BD",x"F5",x"7E",x"96",x"77",x"27",x"11",x"E6",x"67",
    x"85",x"41",x"26",x"29",x"8D",x"58",x"E4",x"84",x"27",x"02",x"C6",x"01",x"5A",x"20",x"1B",x"BD",
    x"F7",x"ED",x"E6",x"67",x"8D",x"4C",x"1F",x"98",x"E6",x"84",x"7C",x"A7",x"C0",x"A4",x"84",x"26",
    x"05",x"C4",x"0F",x"53",x"20",x"04",x"54",x"54",x"54",x"54",x"E7",x"64",x"39",x"44",x"25",x"0D",
    x"54",x"E6",x"84",x"25",x"04",x"54",x"54",x"54",x"54",x"C4",x"0F",x"20",x"ED",x"BD",x"F7",x"E4",
    x"BD",x"F5",x"52",x"4F",x"E5",x"84",x"27",x"02",x"86",x"02",x"7A",x"A7",x"C0",x"E5",x"84",x"27",
    x"01",x"4C",x"1F",x"89",x"20",x"D4",x"96",x"77",x"85",x"40",x"26",x"22",x"D6",x"33",x"85",x"20",
    x"26",x"08",x"CE",x"F6",x"61",x"C4",x"07",x"E6",x"C5",x"39",x"CE",x"F6",x"61",x"C4",x"03",x"E6",
    x"C5",x"96",x"79",x"84",x"03",x"85",x"01",x"27",x"04",x"54",x"54",x"54",x"54",x"39",x"EC",x"65",
    x"54",x"D6",x"29",x"25",x"06",x"58",x"58",x"58",x"58",x"4F",x"39",x"C4",x"0F",x"39",x"96",x"77",
    x"85",x"60",x"26",x"1F",x"1F",x"20",x"86",x"28",x"3D",x"1E",x"01",x"44",x"56",x"44",x"56",x"54",
    x"0D",x"77",x"2A",x"0C",x"54",x"30",x"8B",x"BD",x"F7",x"E4",x"24",x"03",x"7A",x"A7",x"C0",x"39",
    x"30",x"8B",x"39",x"1F",x"20",x"86",x"28",x"3D",x"1E",x"01",x"34",x"04",x"54",x"54",x"30",x"8B",
    x"BD",x"F7",x"E4",x"96",x"77",x"85",x"20",x"27",x"0E",x"96",x"79",x"85",x"02",x"27",x"03",x"7A",
    x"A7",x"C0",x"35",x"04",x"7E",x"F5",x"9F",x"86",x"04",x"3D",x"E0",x"E0",x"53",x"5C",x"54",x"54",
    x"20",x"C8",x"BD",x"F7",x"D0",x"96",x"29",x"2B",x"12",x"EA",x"84",x"E7",x"84",x"D6",x"19",x"C5",
    x"10",x"26",x"23",x"48",x"48",x"48",x"48",x"C6",x"0F",x"20",x"10",x"53",x"E4",x"84",x"E7",x"84",
    x"D6",x"19",x"C5",x"10",x"26",x"10",x"43",x"84",x"0F",x"C6",x"F0",x"7A",x"A7",x"C0",x"E4",x"84",
    x"E7",x"84",x"AB",x"84",x"A7",x"84",x"39",x"96",x"77",x"85",x"40",x"10",x"26",x"00",x"42",x"85",
    x"20",x"10",x"26",x"FF",x"C0",x"44",x"24",x"BA",x"BD",x"F7",x"E4",x"96",x"29",x"84",x"03",x"44",
    x"1F",x"98",x"26",x"10",x"25",x"0E",x"53",x"E4",x"84",x"E7",x"84",x"43",x"7A",x"A7",x"C0",x"A4",
    x"84",x"A7",x"84",x"39",x"25",x"06",x"EA",x"84",x"E7",x"84",x"20",x"EF",x"26",x"07",x"53",x"E4",
    x"84",x"E7",x"84",x"20",x"04",x"EA",x"84",x"E7",x"84",x"7A",x"A7",x"C0",x"AA",x"84",x"A7",x"84",
    x"39",x"24",x"03",x"86",x"F0",x"8C",x"86",x"0F",x"A4",x"84",x"A7",x"84",x"EA",x"84",x"E7",x"84",
    x"39",x"80",x"40",x"20",x"10",x"08",x"04",x"02",x"01",x"34",x"7E",x"86",x"20",x"1F",x"8B",x"CC",
    x"01",x"01",x"34",x"06",x"4F",x"E6",x"68",x"D0",x"35",x"22",x"0E",x"26",x"09",x"0D",x"36",x"26",
    x"05",x"35",x"06",x"7E",x"F6",x"F4",x"60",x"61",x"50",x"DD",x"46",x"EC",x"65",x"93",x"32",x"22",
    x"07",x"60",x"E4",x"43",x"53",x"C3",x"00",x"01",x"DD",x"44",x"9E",x"32",x"10",x"9E",x"34",x"10",
    x"93",x"46",x"22",x"28",x"D6",x"47",x"27",x"48",x"54",x"50",x"86",x"FF",x"31",x"21",x"6D",x"61",
    x"2A",x"02",x"31",x"3E",x"D3",x"44",x"2B",x"0A",x"30",x"01",x"6D",x"E4",x"2A",x"02",x"30",x"1E",
    x"93",x"46",x"BD",x"F4",x"A3",x"10",x"AC",x"67",x"27",x"26",x"20",x"E0",x"43",x"53",x"C3",x"00",
    x"01",x"47",x"56",x"30",x"01",x"6D",x"E4",x"2A",x"02",x"30",x"1E",x"D3",x"46",x"2B",x"0A",x"31",
    x"21",x"6D",x"61",x"2A",x"02",x"31",x"3E",x"93",x"44",x"BD",x"F4",x"A3",x"AC",x"65",x"26",x"E3",
    x"32",x"62",x"35",x"FE",x"9C",x"32",x"22",x"08",x"27",x"5B",x"DE",x"32",x"1E",x"13",x"DF",x"32",
    x"34",x"10",x"96",x"77",x"85",x"60",x"26",x"5E",x"DC",x"32",x"44",x"56",x"44",x"56",x"54",x"34",
    x"04",x"1F",x"10",x"44",x"56",x"44",x"56",x"54",x"E0",x"E0",x"27",x"3B",x"34",x"04",x"9E",x"32",
    x"BD",x"F5",x"7E",x"BD",x"F5",x"46",x"58",x"5A",x"BD",x"F6",x"07",x"0D",x"77",x"2A",x"0E",x"B6",
    x"A7",x"C0",x"44",x"24",x"05",x"7A",x"A7",x"C0",x"20",x"05",x"7C",x"A7",x"C0",x"30",x"01",x"C6",
    x"FF",x"6A",x"E4",x"2E",x"E3",x"35",x"04",x"EC",x"E1",x"BD",x"F5",x"55",x"5A",x"53",x"BD",x"F6",
    x"07",x"AE",x"63",x"9F",x"32",x"35",x"FE",x"9E",x"32",x"BD",x"F4",x"A3",x"30",x"01",x"AC",x"E4",
    x"2F",x"F7",x"32",x"62",x"20",x"EB",x"DC",x"32",x"54",x"54",x"34",x"04",x"1F",x"10",x"54",x"54",
    x"E0",x"E0",x"27",x"E3",x"34",x"04",x"9E",x"32",x"8D",x"31",x"6A",x"E4",x"2F",x"1F",x"BD",x"F5",
    x"7E",x"96",x"77",x"85",x"20",x"26",x"33",x"D6",x"29",x"58",x"58",x"58",x"58",x"DA",x"29",x"E7",
    x"84",x"7A",x"A7",x"C0",x"E7",x"80",x"7C",x"A7",x"C0",x"6A",x"E4",x"2E",x"F2",x"35",x"04",x"EC",
    x"E4",x"C4",x"FC",x"1F",x"01",x"EC",x"E1",x"8D",x"05",x"20",x"A6",x"1F",x"10",x"53",x"C4",x"03",
    x"5C",x"BD",x"F4",x"A3",x"30",x"01",x"5A",x"26",x"F8",x"39",x"C6",x"F0",x"BD",x"F5",x"61",x"34",
    x"04",x"E6",x"E4",x"BD",x"F6",x"07",x"30",x"01",x"6A",x"61",x"2E",x"F5",x"35",x"04",x"20",x"CD",
    x"96",x"77",x"2B",x"18",x"27",x"0E",x"85",x"02",x"26",x"19",x"85",x"04",x"26",x"06",x"96",x"79",
    x"84",x"01",x"26",x"0F",x"B6",x"A7",x"C0",x"8A",x"01",x"B7",x"A7",x"C0",x"39",x"96",x"79",x"84",
    x"01",x"26",x"F1",x"B6",x"A7",x"C0",x"84",x"FE",x"20",x"EF",x"0D",x"79",x"10",x"2B",x"04",x"E2",
    x"A6",x"C4",x"84",x"02",x"34",x"02",x"BE",x"EF",x"F4",x"8C",x"58",x"12",x"26",x"05",x"86",x"02",
    x"B7",x"21",x"94",x"8E",x"04",x"E1",x"BD",x"F4",x"75",x"A6",x"C4",x"84",x"02",x"A1",x"E0",x"26",
    x"D9",x"8B",x"FF",x"39",x"0D",x"79",x"10",x"2B",x"04",x"CD",x"1A",x"50",x"9E",x"67",x"34",x"18",
    x"8E",x"F9",x"3B",x"9F",x"67",x"86",x"A7",x"1F",x"8B",x"10",x"8E",x"20",x"CD",x"8E",x"03",x"70",
    x"86",x"FF",x"D6",x"E7",x"2A",x"FC",x"D6",x"E7",x"2B",x"FC",x"A7",x"42",x"BD",x"F4",x"75",x"6D",
    x"C4",x"8E",x"06",x"49",x"86",x"01",x"97",x"E4",x"96",x"E5",x"1C",x"BF",x"BD",x"F4",x"75",x"1A",
    x"40",x"CE",x"A7",x"C0",x"1C",x"EF",x"86",x"FE",x"A7",x"42",x"0F",x"E4",x"35",x"08",x"10",x"8C",
    x"20",x"D0",x"23",x"77",x"1F",x"23",x"A6",x"5E",x"80",x"06",x"A8",x"5E",x"84",x"07",x"A8",x"5E",
    x"A7",x"5E",x"AE",x"5D",x"86",x"80",x"A5",x"C2",x"27",x"14",x"44",x"A5",x"C4",x"26",x"0F",x"A6",
    x"5F",x"84",x"38",x"81",x"20",x"25",x"07",x"81",x"38",x"26",x"50",x"30",x"88",x"C0",x"AF",x"C3",
    x"11",x"83",x"20",x"CD",x"26",x"D0",x"4F",x"D6",x"78",x"DD",x"44",x"31",x"3D",x"5F",x"AE",x"C1",
    x"A6",x"C0",x"30",x"89",x"01",x"40",x"AC",x"C4",x"22",x"37",x"30",x"08",x"AC",x"C4",x"25",x"31",
    x"30",x"18",x"AF",x"C4",x"A7",x"42",x"5C",x"20",x"2B",x"6A",x"6B",x"30",x"89",x"01",x"40",x"1F",
    x"10",x"93",x"44",x"2B",x"0A",x"10",x"83",x"01",x"40",x"25",x"06",x"CC",x"01",x"3F",x"8C",x"DC",
    x"27",x"0D",x"77",x"2A",x"02",x"58",x"49",x"ED",x"68",x"4F",x"21",x"43",x"35",x"10",x"9F",x"67",
    x"39",x"5D",x"26",x"0A",x"34",x"40",x"10",x"AC",x"E1",x"26",x"B3",x"5D",x"27",x"ED",x"86",x"03",
    x"3D",x"50",x"33",x"C5",x"EC",x"C4",x"10",x"83",x"FA",x"00",x"24",x"DF",x"8E",x"FF",x"F5",x"30",
    x"0A",x"83",x"0C",x"80",x"24",x"F9",x"C3",x"0C",x"80",x"30",x"01",x"83",x"01",x"40",x"24",x"F9",
    x"C3",x"01",x"40",x"AF",x"6A",x"1F",x"01",x"E6",x"42",x"C5",x"80",x"27",x"A2",x"8C",x"00",x"3F",
    x"25",x"97",x"8C",x"00",x"FF",x"23",x"98",x"6C",x"6B",x"20",x"A4",x"0D",x"E5",x"CC",x"F9",x"44",
    x"FD",x"20",x"67",x"3B",x"DE",x"E4",x"10",x"8C",x"20",x"E1",x"24",x"0A",x"DC",x"E6",x"58",x"2A",
    x"05",x"EF",x"A1",x"A7",x"A0",x"3B",x"8E",x"00",x"01",x"3B",x"1A",x"D0",x"96",x"3C",x"D6",x"3A",
    x"34",x"02",x"44",x"44",x"AB",x"E0",x"3D",x"1F",x"02",x"E6",x"64",x"C4",x"0F",x"27",x"0C",x"8E",
    x"F9",x"C4",x"E6",x"85",x"96",x"3F",x"4A",x"26",x"02",x"C0",x"02",x"1F",x"98",x"DD",x"44",x"27",
    x"10",x"9E",x"3E",x"E6",x"41",x"CA",x"01",x"E7",x"41",x"D6",x"45",x"8D",x"20",x"30",x"1F",x"26",
    x"F2",x"9E",x"3E",x"E6",x"41",x"C4",x"FE",x"E7",x"41",x"D6",x"44",x"8D",x"10",x"30",x"1F",x"26",
    x"F2",x"DC",x"44",x"9B",x"3D",x"25",x"EA",x"D0",x"3D",x"22",x"D2",x"20",x"E4",x"D7",x"46",x"5A",
    x"26",x"FD",x"D6",x"46",x"27",x"08",x"DB",x"47",x"D1",x"47",x"D7",x"47",x"24",x"04",x"31",x"3F",
    x"27",x"01",x"39",x"35",x"86",x"B0",x"A5",x"9C",x"92",x"89",x"81",x"78",x"71",x"6A",x"63",x"5D",
    x"57",x"51",x"CE",x"A7",x"CC",x"96",x"42",x"8A",x"D0",x"1F",x"8A",x"25",x"0A",x"29",x"08",x"96",
    x"42",x"97",x"43",x"4F",x"39",x"43",x"39",x"86",x"04",x"95",x"43",x"27",x"F8",x"A6",x"54",x"8A",
    x"04",x"A7",x"54",x"86",x"0A",x"97",x"7E",x"34",x"04",x"EC",x"42",x"84",x"FB",x"C4",x"FB",x"ED",
    x"42",x"CC",x"F3",x"33",x"ED",x"C4",x"EC",x"42",x"8A",x"04",x"CA",x"04",x"ED",x"42",x"35",x"04",
    x"96",x"42",x"85",x"02",x"26",x"18",x"8D",x"74",x"EC",x"42",x"84",x"FB",x"C4",x"FB",x"ED",x"42",
    x"5F",x"4F",x"ED",x"C4",x"EC",x"42",x"8A",x"04",x"CA",x"04",x"ED",x"42",x"4F",x"39",x"3F",x"06",
    x"10",x"9E",x"27",x"0D",x"77",x"2B",x"12",x"C6",x"07",x"8D",x"51",x"E6",x"A0",x"E7",x"C4",x"8D",
    x"57",x"10",x"8C",x"1F",x"40",x"25",x"F4",x"20",x"CF",x"8E",x"FA",x"AF",x"8D",x"1F",x"86",x"28",
    x"8D",x"20",x"6A",x"54",x"8D",x"1C",x"6C",x"54",x"31",x"21",x"4A",x"26",x"F3",x"31",x"A9",x"01",
    x"18",x"10",x"8C",x"1F",x"40",x"25",x"E2",x"8D",x"04",x"20",x"AD",x"8D",x"1F",x"E6",x"80",x"26",
    x"FA",x"39",x"C6",x"08",x"34",x"26",x"C6",x"80",x"68",x"A4",x"24",x"02",x"6C",x"A4",x"56",x"31",
    x"A8",x"28",x"24",x"F4",x"8D",x"06",x"35",x"26",x"5A",x"26",x"E9",x"39",x"34",x"04",x"E7",x"C4",
    x"E8",x"C4",x"C4",x"03",x"35",x"04",x"26",x"F4",x"58",x"58",x"CA",x"03",x"E7",x"41",x"A6",x"43",
    x"88",x"08",x"A7",x"43",x"88",x"08",x"A7",x"43",x"A6",x"43",x"2A",x"FC",x"6D",x"41",x"39",x"0A",
    x"1B",x"39",x"1B",x"46",x"31",x"36",x"30",x"1B",x"47",x"36",x"34",x"30",x"00",x"0A",x"1B",x"36",
    x"00",x"E6",x"4C",x"4D",x"27",x"06",x"86",x"40",x"54",x"54",x"54",x"54",x"C4",x"0F",x"8E",x"FA",
    x"D7",x"E6",x"85",x"E7",x"64",x"8B",x"40",x"A4",x"4D",x"81",x"01",x"39",x"04",x"02",x"03",x"00",
    x"06",x"08",x"07",x"00",x"05",x"01",x"00",x"86",x"A7",x"1F",x"8B",x"10",x"8E",x"20",x"82",x"A6",
    x"A4",x"1F",x"8A",x"25",x"1C",x"29",x"1A",x"27",x"0E",x"86",x"10",x"A7",x"21",x"96",x"EA",x"8A",
    x"02",x"97",x"EA",x"96",x"E9",x"20",x"12",x"86",x"04",x"A5",x"21",x"26",x"12",x"A7",x"21",x"20",
    x"10",x"86",x"04",x"A5",x"21",x"27",x"08",x"8D",x"45",x"4F",x"39",x"86",x"80",x"A7",x"21",x"43",
    x"39",x"1A",x"10",x"4F",x"E6",x"23",x"1F",x"03",x"A6",x"22",x"84",x"E1",x"88",x"61",x"8B",x"40",
    x"1C",x"FE",x"46",x"24",x"02",x"8A",x"80",x"33",x"C6",x"1F",x"30",x"D7",x"EB",x"E6",x"22",x"C4",
    x"1C",x"58",x"58",x"58",x"96",x"EA",x"84",x"10",x"8A",x"09",x"34",x"02",x"EA",x"E0",x"D7",x"EA",
    x"53",x"D8",x"EA",x"5C",x"26",x"C5",x"CE",x"F1",x"84",x"FF",x"20",x"64",x"20",x"BB",x"A6",x"A4",
    x"85",x"02",x"26",x"11",x"96",x"E9",x"85",x"10",x"27",x"FA",x"86",x"3C",x"4A",x"96",x"E9",x"48",
    x"2B",x"F2",x"D7",x"E8",x"39",x"96",x"E9",x"85",x"08",x"26",x"15",x"1A",x"10",x"E6",x"22",x"54",
    x"54",x"25",x"03",x"48",x"2B",x"06",x"96",x"EA",x"8A",x"08",x"97",x"EA",x"32",x"62",x"20",x"8F",
    x"D6",x"E8",x"84",x"03",x"26",x"E5",x"E7",x"66",x"39",x"0F",x"7F",x"C6",x"08",x"F7",x"A7",x"DD",
    x"8E",x"EF",x"E0",x"E6",x"80",x"27",x"06",x"C1",x"04",x"2D",x"07",x"27",x"15",x"8C",x"EF",x"F4",
    x"26",x"F1",x"4F",x"8E",x"A5",x"5A",x"BC",x"EF",x"FB",x"26",x"01",x"43",x"C6",x"28",x"F7",x"A7",
    x"DD",x"39",x"0C",x"7F",x"5F",x"8D",x"19",x"8E",x"EF",x"E0",x"E6",x"84",x"C1",x"20",x"26",x"04",
    x"30",x"01",x"20",x"F6",x"8D",x"28",x"C6",x"0D",x"3F",x"02",x"C6",x"0A",x"3F",x"02",x"20",x"D2",
    x"34",x"14",x"8E",x"FC",x"51",x"9F",x"70",x"8E",x"FC",x"43",x"8D",x"12",x"C6",x"30",x"EB",x"E0",
    x"3F",x"02",x"C6",x"20",x"3F",x"02",x"35",x"90",x"8D",x"E6",x"20",x"02",x"8D",x"07",x"E6",x"80",
    x"C1",x"04",x"26",x"F8",x"39",x"5D",x"2A",x"39",x"3F",x"06",x"FE",x"20",x"70",x"C0",x"80",x"86",
    x"08",x"3D",x"33",x"CB",x"7F",x"20",x"30",x"10",x"BE",x"20",x"21",x"C6",x"08",x"37",x"02",x"A7",
    x"A4",x"31",x"A8",x"D8",x"5A",x"26",x"F6",x"C6",x"08",x"10",x"BE",x"20",x"21",x"3F",x"04",x"B6",
    x"20",x"2B",x"A7",x"A4",x"31",x"A8",x"D8",x"5A",x"26",x"F8",x"7C",x"20",x"1C",x"7C",x"20",x"22",
    x"39",x"3F",x"82",x"1B",x"44",x"1B",x"53",x"80",x"81",x"81",x"82",x"1B",x"40",x"1B",x"58",x"20",
    x"04",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",
    x"FF",x"C6",x"A7",x"1F",x"9B",x"4D",x"2A",x"21",x"0D",x"E7",x"2A",x"FC",x"0D",x"E7",x"2B",x"FC",
    x"10",x"8E",x"02",x"00",x"31",x"3F",x"26",x"FC",x"0F",x"DB",x"10",x"8E",x"00",x"10",x"EC",x"81",
    x"D7",x"DA",x"97",x"DA",x"31",x"3F",x"26",x"F6",x"39",x"48",x"34",x"02",x"8D",x"29",x"C6",x"0A",
    x"5A",x"26",x"FD",x"12",x"A6",x"E4",x"97",x"DB",x"1F",x"10",x"D4",x"DA",x"94",x"DA",x"34",x"06",
    x"1F",x"20",x"AA",x"E0",x"EA",x"E0",x"AC",x"81",x"1F",x"01",x"35",x"02",x"97",x"DB",x"1F",x"10",
    x"D7",x"DA",x"97",x"DA",x"AF",x"66",x"39",x"86",x"20",x"B5",x"A7",x"E7",x"27",x"FB",x"B5",x"A7",
    x"E7",x"26",x"FB",x"5A",x"34",x"7E",x"3D",x"3D",x"1A",x"00",x"35",x"7E",x"B5",x"A7",x"E7",x"27",
    x"F2",x"39",x"B6",x"A7",x"CC",x"84",x"03",x"27",x"0B",x"81",x"02",x"22",x"03",x"27",x"02",x"4F",
    x"39",x"4F",x"43",x"39",x"1A",x"05",x"39",x"96",x"79",x"85",x"40",x"27",x"1C",x"A6",x"4F",x"84",
    x"FB",x"A7",x"4F",x"E6",x"4D",x"C5",x"04",x"34",x"01",x"C4",x"FB",x"E7",x"4D",x"8A",x"04",x"A7",
    x"4F",x"35",x"01",x"27",x"06",x"86",x"1F",x"A7",x"4E",x"43",x"39",x"4F",x"34",x"01",x"1A",x"50",
    x"96",x"77",x"2A",x"08",x"DC",x"7A",x"8D",x"26",x"02",x"7F",x"20",x"12",x"85",x"60",x"27",x"08",
    x"DC",x"7A",x"8D",x"1A",x"00",x"9F",x"20",x"06",x"DC",x"7A",x"8D",x"12",x"01",x"3F",x"DD",x"7A",
    x"ED",x"67",x"DC",x"7C",x"8D",x"08",x"00",x"C7",x"DD",x"7C",x"ED",x"69",x"35",x"81",x"35",x"10",
    x"4D",x"2A",x"02",x"4F",x"5F",x"10",x"A3",x"84",x"23",x"02",x"EC",x"84",x"6E",x"02",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F1",x"D9",
    x"01",x"00",x"F0",x"53",x"F0",x"53",x"F0",x"A1",x"F0",x"B9",x"F0",x"9D",x"F0",x"53",x"F1",x"9F");

END PACKAGE;